BSV1    $k�h� �            �+�FV  ���FV  �+�FV  �+�FV                      �                                                         `	��Z  � $ B   �  Ji BB      �     ��              �X       Ptj      8t j      X       @                �  |�s    |�s                  ��e	���  j/=�0N
��Hm,
��e�%�O�gF��H�!m,��eO��hF� H�!m,��eO��L
�� @�-k%J!��O1�4��gF��` �e	�=�5�5K/=�0M�gF��` N-��B f�$�$` ) 1e5�=�$�c)%J)k-�1�5�9�=B1FRJsN�R�V�Z�^UU���<1!�-�B�df�Ip^0s�|�UU�t��U.W�6�W�8]]_vS`9�{UU�� z5]>�::WCr�-�6�[8U�z�UU�w�f-�-J?�G��j ��R�1�QR  ,��S��f{�z�Uv�~/~�	��5�� ��5�R�yZr�~]5�.^7�_��� ��5�R�yZr�~]5�.^7�_�  � � �    � � h     � � j     � � l     � � n     � �       � � D     � � F     � � �    � � �    � �       � M 
      �       �     � @     � @    � P    � P   � H �     � � �     � �       � �       � �       � � �     � � �     � � �     � � �     � �       � � @     � � B    � �       � �       � �      � �      � �      � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   � � U   X � �    � � h      � � j      � � l      � � n      � �       � c �    � s �    � y       , Y �     < Y �     , i �     < i �     8 h         @     
  B              � �       � �       � � &     � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U    � � U            � � � �     �   =�     � �        �  ���3��h<��j<��l<��n<�� 2��D1��F1���3���#�� "�M
3 �5 �7�@3�@s�P��P�H�8���8�� 2�� 2�� 2��>��>��>��>�� 2��@:��Bz�� 2�� 2��"��"��"��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UUX��3��h0��j0��l0��n0�� 2�c�3�s�#�y ",Y�p<Y�p,i�p<i�p8h 2@p
B0 2�� 1�� 1��&1��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ                                �         ��                               UQ  �       ��!     �        ��"    >�~     ~ ��&    �       ~  ��&    �  2    �  ��               �             �  �D                 
�C          Ie`�`��`���Y�� � � �@� @  � �p ��0�0��0p�@�@� �b�"�(��� �. ���O0����������������r g ["��O���f������;?��9y^��� uD�����������������           l            q            ��@            � � �  
        �ۘ�����I~��@�z}        � @   � ��$�DИ�*Sv(L( ?@� � � �$   � � �� � � �`  � � � � � �@� �/�¹�,�g=������D��������_���)�z{��{���`  W���   �j
��0�X�
2�=¶A�0 O �  @ Fb8�x��z��$q��~��}�����s��k�m�	o_� ���А���������-�� 5
` o`�����A���������|��8��^ � �������������ڧ�
���8�gV����@�������������#�#��>B�� ���������                �[?@�3�>������� � 3          ����`$����R�v���p 8 �      	)8<  X@X@t`2 a@`@%��{�������}��{X    @     �                              �����        �   ca�B{d�8�<�٘� � � � � � � �M��-�%B&A�A�!�!� � � � � � � � �d�l�,�k�c٣7*C�C�C�B�� �� � �i�	���ʇ��0�a�  ��_�    `8��g�?     `��g8 �                             �����        �   ca�B{d�8�<�٘� � � � � � � �M��-�%B&A�A�!�!� � � � � � � � �d�l�,�k�c٣7*C�C�C�B�� �� � �i�	���ʇ��0�a�  ��_�    `8��g�?     `��g8 �          �   �          � � 0 �QK�� � KɷT�T�i���?�?����� * �����k?X7U�������V�����                    O=�3\��d]@�	r��?���������"O�1���۵���g�������*�$�J�)�ZF),æ�����7ݱ � ��p�Q���&��ݞ`�8�?�>��w�|%�� � � ���?���A>�v��3�q�ߔK���?�������k���:**f   
!! ! A 4���(6:<�fD�   � � � �|�y�1з@���+�,�� � ���~�p�p��"�"�2�s����� � � � � �   ?�O��єQ�P� � D d d � � � � � j������hd�z�:!>!~|�L#F)p�x�� �AK�����!��� ����Ȑ�(�d��|�8 8 x � � � � � �t�0�(� � 5��@�q��'���?����� WA�G�	^�v�\��������������d(07T}�}��`|��7/k�/��?�?���*.��.�nGg�����������������03
���pt4���{?�����P �ۋ}T�՝��GI�����t���*�jѸ]J�vc���R{h���O����$��3� �g�3���;,���������U�2���p��9�9�1�#h`wg�G�_��� � � ��� ba�yx�@�>����a�a�y	��>�Qn����h�$�&�*_�����;ȹH� ����rd�8"<��  � � ���`� �aqP#Z&\$R"W'u
������� �4{�;�;��� /���q�� � � �  a�e�~���>��`�$�����	�0��"�b�.�	����� � � � � �?  ~��@�A�J!�]��*�&�������_�/��2ݺ�r�������gؿ��� �   �p��R����q �`�������o������=�p��R �zր��?�������������'�Qm   � � ?����Z�������������@[� �� ����~������w�����Q � �@� ��� 4 �������������������][.vQ����~���������������!/H#H<[~/�/� � � ��� ��5���ؚe����� ? �X��=�/�����H�T�W�/�/� p p t�� ��c�3��ޘg�����  ? �X��=��ck6�;�e�b!�`a`� � � ��|����X�[�8�hǊ�\�]�/ , < � � � � 4<>c�b!�`a`���`�ă|����X�Y�(�HƊ�M�M�   ? � � � � ~�_�����@� W�������� � ���/���H��r�:S�~����7�q v6"�����۷�C~������[�*�$�J��VրV� ]O^U���C�����������nѾ\C�˔���ՊՊ�Ω־>~         `8��g�?     `��g8 �          �   �          � � 0 U���l?� �g�? ����o��g8 �\C�˔���ՊՊ�Ω־>~         `8��g�?     `��g8 �          �   �          � � 0 U���l?� �g�? ����o��g8 ��9�,_�o��7���V��� �8�0�� �A�`�>���2��q����������c�����u#N9�M�,ѮL��Np��������S��o�?                             �����        �   �d=�L̹H��aq� C�c�c '@�@�������f��� � � � � � � ���p�?P�x�x�X����8<<<�����%�"��8�0�pLp��x���Z�)�,�6���Z[I1 p p ` a � � � ��
�i� �X~�_	���������������Z�S���Z���޿������?�?�����������             L3F9h�n��2��6����!�!�a�A� � � �hp`| FD0  0 � � � �8�<����]Z�U��{)_�����������������'6����6��������[����������������%UQQ�7��>�f�(���������������o���H�`��F�G���-7?��?~�^�� <'_     > C � 4���(��:;��    � � � �  � � � �@ @  @�@� � � � � � � � &�4ȴI�)����]r���~�� �x�|Z$S�               �$�-�l�Hj�k٫�8� �� ���� ��y�����¿��0�A��y���g�/_0�p   <Br�y��1��xg   <~Q��1��f� �����   � � � x�t�               �$�-�l�Hj�k٫�8� �� ���� ��y�����¿��0�A��y���g�/_0�p   <Br�y��1��xg   <~Q��1��f� �����   � � � x�t�� �����Nn��� �         0Rd}��/Q,�J  < n �   ���<���'�;�r���<�� � øG�o�o��m�-�-�%B6A6���� � � � � ����@� @� ��  � �@�� � � � � � � @�   <Br�y��>�0�   <~Q���n�b�y�Ƴ���G#�y�5��=���4���������;��3h��&���/ 3L��B'�#�/ן����`�`����� v ���f����������A>�?�9�1R!l@?D;� �������<�C�`��@�X��-��� �� ��_���          u0U����@�@� � ��l���� � ��j ~ ��d�z�:�a>��<��b]zEjeAN! ZD�J�J�j�I�	�	�K�����K7����|CmC|�|��    � � 7 >�yt7K?@'U��������� � �	e�%� ��r����\���<����#d��w ���+�,π�?@�o��~�p�p���������?�?�?��� �   @� � � � � �@� �@� � � � � �@�@��M�e�e�nA>@?J4@>�5�5�5�6����z۸1��C����kJw���g�����[�n���ZF),æ�⮲��{�� � ��p�Q�}������`�8�?�>��w��� � � ���?���A>�v�6���K�H�k$��?���[��������`�8�?�>��w�|�� � � ���?���                   �&�G�|����Cy`[B� �`�$�4�̂n�L��4�A�A�A�C�@�@0? ? ? ? ? ? ����a�!�#�#^�����"ݣ\�����r���eb�c  � � ��c�c�aqS#S#X �"� u
��������4�t�d�d[$W(ȷ��q�`�`ߠߠ���_f�f�f�g�c�s�3�� � � � � � � � C<�>�9�1X!bd`� ������� �� � �  � �    @�� � � � �     B<�<�>�n�n�~�n��������}��� � � � ��}�l�P�`����?��R� � ��@��zZ����R� �?������������������������������������������7��� � � � ����6�
���������A>�v��1�y�� K ��?�����������=�=�uk���? ���������?�������%�"��8�0�pLp��x���Z�)�,�6���Z[I1 p p ` a � � � 	5����������}}}�����3h��$��K7@?3L��s$�!�*�L�H��`�@>�>��΁r���.����@ <�C�p<�¨�������� � !    2BRb����� �� �!� � ?  �  � � `�8�8�8�8�}�} ����������$؁~����������������������%�5I5�����������������a�!�#�#^�����"ݣ\�����r���eb�c  � � ��c�c�aqS#S#X �"� u
��������4�t�d�d[$W(ȷ��q�`�`ߠߠ��G?O?O?o?o???����/�/�?�?��$�-�l�Hj�k٫�8� �� ���� ��9�,_�O�N�&ƯO�v��� ��&ٮQ�a�d=�5l�����!� C�C�c � � � ���<�Br�y����vq��9�~�.8���p��h�x�t�7E����X�T�[�X�� � y�t���V���➡�� ? ? ? @@[|StWp70g F��� � � � � � ��������f��� � � � � � � ���p �PoxG���������<< � �����5�>������������������X�<�r��~�v�v���9�>�~�q�b�~P�	5����������}}}�����3h��$��K7@?3L��s$�!�*�L�H��`�@>�>��΁r���.����@ <�C�p<�¨�������� � !    ��R� � ��@��zZ����R� �?���������0��P�@����� נ�����|�|���~���I�J3°Q�H]*Y��#�g�g�n�.�������
4j�t�r�����r]jEjeAN! ZD�Z�J�j�I�	�	�K��	�	��I5����|CmC~�~��    � � w@~����K?@'U������������� �	E�e���s����\���<����#d&�6ȷH�o�p ������?�?�?�q�p�\CTK�U�U�1N)V���� � � � � ��7��� � � � ����6�
����������1�a�A��2�3�0�ZR��"�!�!�!�C�c��0�|�~�.��G�����;�~�g�"��?C��������������?�������������^�����������������������������>�~�t��������?��~��D������.���N��������?��N���N���������������������������������������Ƴ��G�9���=�������������{��4�A�A�A�Ü���0? ? ? ? ? ? ����a�!�#�#^�����"ݣ\�����r���eb�c  � � ��c�c�aqS#S#X �"� u
��������4�t�d�d[$W(ȷ��1�q�`�`ߠߠ�?��_f�f�b�s�u�U��� � � � � � � � A>�?�9�1R!l@?D;� ��������x�
��)�+�uľ�����������������X�p�p�Q���vc�������� ����{�7�wg?C��C�S������������������������������������}��� � � � ��}�l�P�`����?���������������������������������������������������������������������������������������������������"O�1� ����kHg���������{�o���ZF),æ���_� � � ��p�Q�������	5�	����?�<� �}}}�������� �/�ow�[S������������� � �����%����������  *�L�G��L�g�3dX�� � � �����������#2u��T2a���&��Џ� �?�� �0� � � ���[S������������� �  �� � ��%����������  *�L�G�*��C�� �� � � ����������T32���T3`���  ��   �?��� �. ��=Q�P���������������r g;�4L%��?0���������G�k��Ϡ 2*z�X�e�3$^����́�����������@Q�#d��).:<�����Qu���?��                         ���Hy 3 �       G � � ,      0 `ag����Rs      � � h j �            � �                �    	n7� <    & b g x q�$�1�B��vf2 � � 9 y | � � jـB��$j & �V"L� o 1 � � � � �  ����&Lt`��t�p � 0  � �  2 16`O ?x�$�]/�?�H   � � � " o ,ek���M��!�0� �  � " 6 ^ � � ��2�����2�8� < , & � t L � 
&�28 � �X�c��8� � � � � s K G �~&)    � � f  ?     ����A?,����KO j � � # � � ? �}�z��4�:m�A� �D , > K � m � � ��`�tH4< �`    � � � � � � �   �� �/�ow�[S������������� � �����%����������  *�L�G��L�g�3dX�� � � �����������#2u��T2a���&��Џ� �?�� �0� � � ���[S������������� �  �� � ��%����������  *�L�G�*��C�� �� � � ����������T32���T3`���  ��   �?��� �. ��=Q�P���������������r g;�4L%��?0���������G�k��Ϡ 2*z�X�e�3$^����́�����������@Q�#d��).:<�����Qu���?��                         ���Hy =�       G � �"     0 `ag����f      � � h b�<           � �                �                          ���Hy =�       G � �"     0 `ag����f      � � h b�<           � �                � o7� <  & b g x }�$�1�B��{9vf2� � 9 I0x�0�zـB��$m#�V"��o 1 � ���1� �܈��&Lt`��t�p  �0� � �  2 16`L;�'�]/�?�H  }��� " o -ek���M��!�0�� � " 6 ^ � ]���2�����:�83�<�, &� t D8�8
&�2�������c��8� � ��'�s K G �~&)    � � f  ?     ����A?,����KO j � � # � � ? ��}�z��4�:m�A� �D, > K � m � � ��`�tH4< �`    � � � � � � �   ��gV�۸�s�RS���������������������d�By�Ҫ���w}���߽���(�`*�L�G��L�g�3dX�� � � �����������#2u��T2a���&��Џ� �?���^!�a7F.N�mo�����ƹ̱���ꑃ8d�lb��t�x������c���7���O&F�B@=J��[wZͰƹ½����=������d��YF�	�]����'�dE��������� �|�z�v�n�^�>� �  ||zzvvnn^^>>   �|�z�v�n�^�>� �  ||zzvvnn^^>>   �|�z�v�n�^�>� �  ||zzvvnn^^>>   �|�z�v�n�^�>� �  ||zzvvnn^^>>  #̤@S��Y�B��K�� �<�l�d�$�8 ; ~1�&�hg�@�� ��N � �p`�G��p�  �Pئ�� �_��@� � I D�|�td8� ��FW��2�0Ýb�g ��l�L�N�<� � �&�9`�)��S"����y � � � � � I              (,                       �  9          �          @ q 3           D   �  4 ! ��                     
                    ��L�f�`Mb_     & d   ~1�6�s���,J�� ��N � � < � J �  ��D�� |����7 � � � Y �   �G7l��@�&~�� � � r >  � d ��ʀ2�x��B9�"�| } % ' } � � �               ��ҍ�V�r�0� r " b � � � � �  X�%�B�@��vQ.�� � � � � � � � ��F{��:�V�b�g � � � � � � � N �`��3����%� �   < � � �                                  !,�@��      D ' ܬ��s��7  ~a#  � �  � � �  �P>o��� � �< � � r >  � � @;p@��� B9�3�"� �  '  � � �             N1i�7����<���N 	 � | � � � ; ��� �q� ���� � � � � � A O ��3���b������ � � ~  ? � � �|�2_��0�&�j� � � 8 � � � � �@����p�0��@� � I x � � E % � qi��_����  � �  u � � �   �x�9V#� j � �  U �   }n"��D�{�yJ!� � � � � ? � � �o�I�0)X ���8�� � � � � � o  #̬P;ǻi�b��K�� � � � � �  ; �șf�� ���_�� 7   � g b  � ��f� ��z��`~,�� � � N >  � � �z�h��9      � � � �  ! b   N���ÖA��("( 3 s � � w �   	          �@�������Ѐ��@��� ` ` 0   p 8 x n��}�=?;�� � � � � � � � ����j����=-�8{  �   @ @  � ��������) ��F�    _ � { ? � � X�� ���� � � � � � � � ����������) ��F�    _ � { ? ��Y ������ � � � � � � � �����ۏ��G��� ` ` 0   p 8 x ����h����=-�8;  �   @ @ P �  
         ^��}�sꪪ�i�h���     A     #̤@S��Y�B��K�� �<�l�d�$�8 ; ~1�&�hg�@�� ��N � �p`�G��p�  �Pئ�� �_��@� � I D�|�td8� ��FW��2�0Ýb�g ��l�L�N�<� �  � � �� ��o1�� � � � � � � � S�_.`���O�w�@O?������������on}�k�jHw
�ʵ������������������|�?�5����4� � ��8�0��� ~�<B�A��9e���� � � � � � �  �P��w�(�8ǒe� � � � � � � � H�H��Y+�5����B?� � ���������G���M����f�F�+� �`�������������o�*d^�3�.~�'4/����������������W�cH���4�xi�I��� ?��0�������z��<�X&!���6h� � � 7 � �0���`�Cia�Q�:�
m�#���`�`� � � � �  � � �� ��o1�� � � � � � � � S�_.`���O�w�@O?������������on}�k�jHw
�ʵ������������������|�?�5����4� � ��8�0��� ~�<B�A��9e���� � � � � � �  �P��w�(�8ǒe� � � � � � � � H�H��Y+�5����B?� � ���������G���M����f�F�+� �`�������������o�*d^�3�.~�'4/����������������W�cH���4�xi�I��� ?��0�������z��<�X&!���6h� � � 7 � �0���`�Cia�Q�:�
m�#���`�`� � � � � V�H�G@��F�j�[�� � � � � � � � ѭ�%T��5 �I�#P�r � ~ �� �� ʾ�<�o���Z�}y_���������X�~��������fx����������������O�Q��R;G�ik������������������?���}��u�@����V��������@���%�x�q`f���qg����� � �  }`�`����l�\&:��v��0?8<>`�`t88xxૐo�}Bm5+�V$�� ? � � } � � ~ <ìB��Cr��c	��� � � � � � �D	�A��X�}�?��?�����������?�i�|���v�����H�}�m�?�������������_;R�� � j�����������������=�]��Kj�O��p��������������j�.�P���*��o�+@�����������������d��u�������H�����?������������쇪U/�3/;O������� � � � �  �|�z�v�n�^�>� �  ||zzvvnn^^>>   �|�z�v�n�^�>� �  ||zzvvnn^^>>  r��Z�R�@|&����������������������EZ։-H�;����������������?���������@�C���������������v�Y � �Do �������������������=� �h�������-�� � � �`�������� �|�z�v�n�^�>� �  ||zzvvnn^^>>  .z��w5�������� � � }��J ���A��=�=� � � �����o�7��<r,�^d>����������������������J���-������������~�~�~���?��������~@�C����������������A>p?ċ�T����������{�;�����q�#���-_7�7�:-���������o�����F\M�� �H���m�8������B�M�e�������G������?�T��� l�������_����g��u��������������?������k�_�r_��?�?e�	=�����������������\M���j�j�@��H�����O������������G?�}�.����� ������������� �. ��: � v ����������������R g ��� L ��. ������������{����$���T�����i�����������������e � {��@�H���� � � � � � _ � Yۑ�%�Z[,n���j{$ J B � � $ B � d}��dm����T|Z[���  � I % � � A ��R��������F�@I
  R   B ) � Yۑ�/�_O?}���op$ J F � � / F � d}��dm�>�^�~J[���  � A !  � A ��}��C�c�̊5� �0�0� � ��� �<�4�K�$�� � � � � � � � d}��de����N�XY���  � S 3  � a ��%M��_?��y�M}[ � 
 � 
  � � ��Z�=��߾֝�F�@I
  Z   B ) �                                 	          �@�������Ѐ��@��� ` ` 0   p 8 x                                 n��}�=?;�� � � � � � � � ����j����=-�8{  �   @ @  � ��������) ��F�    _ � { ? � � X�� ���� � � � � � � � ����������) ��F�    _ � { ? ��Y ������ � � � � � � � �����ۏ��G��� ` ` 0   p 8 x ����h����=-�8;  �   @ @ P �  
         ^��}�sꪪ�i�h���     A     �C�`������Zx��>      �          �@@�� �   @ � � � � � �                         	=����k�j��s�o$ @ @          ( ( ������������� � | | > > >                                  G##SPj(  � � � o w ~ ?  ZkZ+Z{�s�8J � � � � � � � � ��������/ ߀ �    �  � � �@�D�D� � � `�� � � � � � � � � ��������/!^ > �    � � � � �S�%C�B���o� � � � 0       )!-!������������� � ~  ? ? ?  ZkZkZ{6r  � � � � � � � � � � � UV��Uo��/;O   ( d � D � � �o�o�~�^������ͭ            ix(8�8M�e�'^uLgއ � �   � �    ` ��p 0 � �� � � p � � � � � �d��u�������H�����?������������쇪U/�3/;O������� � � � �  �|�z�v�n�^�>� �  ||zzvvnn^^>>   �|�z�v�n�^�>� �  ||zzvvnn^^>>  r��Z�R�@|&����������������������EZ։-H�;����������������?���������@�C���������������v�Y � �Do �������������������=� �h�������-�� � � �`�������� �|�z�v�n�^�>� �  ||zzvvnn^^>>  .z��w5�������� � � }��J ���A��=�=� � � �����o�7��<r,�^d>����������������������J���-������������~�~�~���?��������~@�C����������������A>p?ċ�T����������{�;�����q�#���-_7�7�:-���������o�����F\M�� �H���m�8������B�M�e�������G������?�T��� l�������_����g��u��������������?������k�_�r_��?�?e�	=�����������������\M���j�j�@��H�����O������������G?�}�.����� ������������� �. ��: � v ����������������R g ��� L ��. ������������{����$���T�����i�����������������e � {��@�H���� � � � � � _ � Yۑ�%�Z[,n���j{$ J B � � $ B � d}��dm����T|Z[���  � I % � � A ��R��������F�@I
  R   B ) � Yۑ�/�_O?}���op$ J F � � / F � d}��dm�>�^�~J[���  � A !  � A � �. ��: � v ����������������R g ��� L ��. ������������{����$���T�����i�����������������e � {��@�H���� � � � � � _ � Yۑ�%�Z[,n���j{$ J B � � $ B � d}��dm����T|Z[���  � I % � � A ��R��������F�@I
  R   B ) � Yۑ�/�_O?}���op$ J F � � / F � d}��dm�>�^�~J[���  � A !  � A ��}��C�c�̊5� �0�0� � ��� �<�4�K�$�� � � � � � � � d}��de����N�XY���  � S 3  � a ��%M��_?��y�M}[ � 
 � 
  � � ��Z�=��߾֝�F�@I
  Z   B ) � q�!q 6A2A�a�`�� � ����� � s�!^!�!bB1@;)ԥ ���� � � � � _kH�� � u�����������������m � ��� U^ � ����������������	���[���y����~�����������������~�{3�+͍��{� � � � � r � � ��%m��M]��i�m}[ �  �   � � � �-��;�#R����������������aZ��� =���3�Y����k�����U��ئ���QO@b�ykT�]ߛ������?���+��dD݀�HT � oD��Ӏ^�������߻�oo=�L,��3�*����� � � � � �@�@� I�8LKS�Ӷ����� � �@� < x  �NZ�	��h���RU� �"��C o � j��i��	(��9������ � { � 3 ss �U�['v9��P�=�� �_������������HDڗ������ � �Z%�Y�w���������t��������� � ���i�w���������� �-��;�#R����������������aZ��� =���3�Y����k�����U��ئ���QO@b�ykT�]ߛ������?���+��dD݀�HT � oD��Ӏ^�������߻�oo=�L,��3�*����� � � � � �@�@� I�8LKS�Ӷ����� � �@� < x  �NZ�	��h���RU� �"��C o � j��i��	(��9������ � { � 3 ss �U�['v9��P�=�� �_������������HDڗ������ � �Z%�Y�w���������t��������� � ���i�w����������� ��d�8@� �������߿������0�p�x�c�}�y��G�� � �� �� i&k�����㔭��%ޞ ��  Z�T&������j�ޖXR � q q # ! ! # ���#���cB{�K��[[ Y q��! 0! �-Catn�)���i����֑�����^Җ�Y�e���7���?��(i�LR@"@b2  Hc���� �@�l��@І �����������SuS�����O��𵄊UWK�_bF{3� �. �	�H2� v�������������ǃ�r g 3Jz�� Y�[�7L�������û �. ��: �w����������������R f�?�{?�u��.Q��������       � �N�	��(�(�r���/?R g ��� L ��z����������������D?�8���M���������������j.G g��[��ڴJ�I�����  �ǚ�7(�N���	8�p���������������H�L��� �������cg*{	���=A��������~���������*�Ʒ+݅�Q��4�����3�{�������� �. �	�H2� v�������������ǃ�r g 3Jz�� Y�[�7L�������û �. ��: �w����������������R f�?�{?�u��.Q��������       � �N�	��(�(�r���/?R g ��� L ��z����������������D?�8���M���������������j.G g��[��ڴJ�I�����  �ǚ�7(�N���	8�p���������������H�L��� �������cg*{	���=A��������~���������*�Ʒ+݅�Q��4�����3�{���������6*t�e�j�������������s���:�p�gi�ؖ\�N[��b}���k�i�����K���� � h&�9�xd�v��������������]�r g�b�l�|؏�0�����������[����9D$�� �	uD�����Ã����������H� ]��0��>�� ����_���!^hK���Ul�D�������������ǃ�;įP� m�g�<�d@�            � ��D�Hs�3���Q�ړ�%O�M�S,5L
��wv"����W��������0_ Gx���fG� �����������������{�v1��,�    �  AG����hQ�� � �^ `���������������c���Oн2� 5 /������������W��-&�\������W���������p�Avz�l�`M���`y���������?�����;3' ����7W����������������CB}�������e��� � @       � @�[Ff�Mzmp��� �������������� M���>�s� ��L�%�(�\��� � � � ;3' ����7W����������������CB}�������e��� � @       � @�[Ff�Mzmp��� �������������� M���>�s� ��L�%�(�\��� � � � ~U��9k�6:)����!� � � � � �T���A� �a ����9�A� � � � g *�;T�0Tt1|`����������������� � \Q~G��1�� � ������pw ߠ��b�� � j ��_�=������������	a��"�����r?�_���l��������(u0hX:�$+Hen8�?�?�_��/�_��?GDl�Ԅ�yA_ObC67����+�?���������7����K�3�#�����    2 �����, M��x�(��{�?����W���/~~�d���5^�KA� �p��%���������������������|����        � �?��������D�Xt���Jvy8; '   � {��4(�8�E�Ԁ������������� ��
5 �I;�m�� � � ��	��O��@� �L҇������ � y�-�I�w��������S*bP���� � �������o���b� l�D҇�)��� � � o�-�I�w����������������A��sc��?�_���Q������<~��(�8n���?�g�?�?��|�
�? � / � ������������������``	Sc�ǲc'u������М�8������ �0���0�T���?�?�?O?�?�_���)���\�\��	_2?��w�I�-�}��� � �)���T�L��WP����w�I�-�}���  ��P*bS�� F\��o�������u��x�8`�	L�T����� � �y�-���������ll� L�S*bP�� � � m�������o��)���\�\��	_2?��w�I�-�}��� � �)���T�L��WP����w�I�-�}���  ��P*bS�� F\��o�������u��x�8`�	L�T����� � �y�-���������ll� L�S*bP�� � � m�������o���~~�	L�T҇�)�� � �y�-�I�w����o��u��똼����zt��  
  C   � k�>�#`�P� �    �  � � � � +/�� � � p�z�� � � � � � � � "b��� � �rra�  � � � � � � KO!�]�  �а � � � � � � / ����������Ԅ1< 7  ?   { � � ��P@Q!������ 6� � � � ~ ? | � ����lt��0���Վ�< 9 � ?   + A CB}�������e�?� � @       � � / _ @ Q����� � � � � � � � ������ܧ������                ^�-��}�~��]<��         �����f���$��88 (p``��mP\�!A1A��燾�? � ? � �  x ` ~�����_�,�d}uu�q [ o   � � ������������|� ��        � �  ��������p ��T@?    � � � � zt�������u����o�   C  
   ��po� x ���׮���� � � �  (   B ��nl�  ���׮��� � � � Q (   C ��~~����u���6� � � � G 
  A ����+p�#:�	��w�Q��� ��������൶��� ��Ed$$�I� D    �F� � ��8����ta \ܲE;�J��	��
� @�y� n�i��
� �����x�
5�&���� ����v� ��> I� ��U��������+p�#:�	��w�Q��� ��������൶��� ��Ed$$�I� D    �F� � ��8����ta \ܲE;�J��	��
� @�y� n�i��
� �����x�
5�&���� ����v� ��> I� ��U����u ��|o�O ��[�aD�  � � � m> ����C3$���\dIr��������π����H��]V�D�z��=�����������c�E�F�aPcOw�`�~����������w���������=  c f � �� (�% J�I��t��������g��?��� � ]��� ��� � � � � � � � ���� �	u��?�5�M � � � � � � � � O�_���
O�_��� ���H ������H �� H������H�����       �      u ������ ������   �  � O�_���
�M� �� ���H(�����ߠ�� H��D��??  �,�      �� � � � u ����>� 88 ���   '����  � � � � � � � �� � � � � � � � &�� ����J�%�������?�o��&4gDw,�X3�u7����������И���.��b]���Dw����Mv�猀����������I�h�+(�g�e:GDs���� ����Pa&����m�M�����w99~������ړ���$ ��   % l n � v   5^�#���   : a � � � � �"��G�1�1��M�� � � � � � � � �\�rG��_��V��#       �@ @ @�@@ ����� � � � � p x ����DC���L�m���O � ? � � � / / S�,pW~���uD�����������������  5^�#���   : a � � � � �"��G�1�1��M�� � � � � � � � �\�rG��_��V��#       �@ @ @�@@ ����� � � � � p x ����DC���L�m���O � ? � � � / / S�,pW~���uD�����������������        y�E         | �       �  �����      � �>                  �              � ��5�� _/�7�����������������{�����h�����        ~��8?�]�z�x�sЁCG''' / [FzD;9q1������#�G�����O� ,���Q�@ @ �� ����������� 8�����?�� �� �_��?���:���^ � �'���?������������F�F�W�[�� � � � � � � � g�0��'d�2L�� �� ��Z��������is��'��=П � �>��o�g�1�W�d�2L�� �� ��Z��������)�s��'��=�_ � �>��o�  
%(      80 @>1N�u��G��������@� � `   ��m��擄&U��c�����)�l��%�����m�ކ���DUѨ�����!�l�H$� G � ��m��Ɠ�~��� �����)�l��$��� �{�U�>��DUѨ�� � ����H � G � �!����1�c���� q  N c � 3 � �m�X�<�S�}�[�m�� � � � � � � � JU�;XkzL��WJk�3������C�����e��C�� �r�{�c� � �`�u�� � � r��e�k�k�`��/�{� � � � � � � � ��m��擄&U��c�����)�l��%�����m�ކ���DUѨ�����!�l�H$� G � ��m��Ɠ�~��� �����)�l��$��� �{�U�>��DUѨ�� � ����H � G � �!����1�c���� q  N c � 3 � �m�X�<�S�}�[�m�� � � � � � � � JU�;XkzL��WJk�3������C�����e��C�� �r�{�c� � �`�u�� � � r��e�k�k�`��/�{� � � � � � � � EV�>\izA��RKc�5�������K������{DY� �&�+�+�� � ����� � � ��1�y�f	{���������������d}��og����H�X[��� �P0�hd};������h鞎� ���	����y�d}��h`���� �L@ڀ� �T/ �? d};-������ )� ����	��x�x�9�� ��c��&O��c��� ������d����{��d@j��� ���� � �� ����`�J���(�� ���� �����<�ÁD���G���	?YA;? ��q�����F���������������yp>8���������D���0O7`YA;?BU�5XkrK��Pm �;������G�����@�*q����}F���>�7���������yp>8� �''�� 2�V����������������� g ����_�� �$� ��?};���� �p�h� ; �A?����������������r G0�z.�7P� ���������������S�����6:d�E�
l�������������t���:�p�g)�ؖT��S��b}���+�a���u�K���`BR��QChE��,+kZڃ���2sv~�׈�A5A�> `�0 
SR4u��44��>��� �''�� 2�V����������������� g ����_�� �$� ��?};���� �p�h� ; �A?����������������r G0�z.�7P� ���������������S�����6:d�E�
l�������������t���:�p�g)�ؖT��S��b}���+�a���u�K���`BR��QChE��,+kZڃ���2sv~�׈�A5A�> `�0 
SR4u��44��>���Q�u�l$�P!�y���������������g ��Q�� � $� �������焄���Z,��/TI ��  ��w���WWKK����"�@!�(B��.#�C�������W��������H �䀰��P P�����̡�x�������2�   SS   ��@  W�� ���    ��)� !1 ���A� $   ��b �9g %%���⪺�����  a@� � �
{G���������������� � �(� �<�>|������� ���}v:D|��8<D�������������������s�5J�\�~	��$�������O��������bf+z��!�%A��������v���������:��f� ;ͅ�Y��4�#���#�{�������)P, 
BRC����@++~~��Dw	{����� 0 �60�: T��DԆ��ڂ���c�Ѐ0�6�P!D�h� ��p��������������*�`@@@     ���� @@@�� B     A@ a`KK  Aa$  � DMb�� ����GGo}���dO���,'>-;%  ` � �   
   ���f����e�M�(_    �   � � � � ���[$��~�{�M�J�     � � � �     "         dO���,'>-;%  ` � �   
   ���f����e�M�(_    �   � � � � ���[$��~�{�M�J�     � � � �     "         q��W�����  |L�  ( � � ! � > � ���(@�P�`�    ��A �    �   �                           ����:?n|3<     � � C  S ?     ��   �         �  � � �       p@(0@hP8 X `x@  ?` `@@`  �͙r��         ���� � � � � �  ��ހ��         (��� � � � � �X@ �� � @       ���� � � � � � �                 � � � � � � � �Ii�@
@   ��9����@� ����     ? H@    0? p@(0@hP8 X `x@  ?` `@@`  �͙r��         ���� � � � � �  ��ހ��         (��� � � � � �X@ �� � @       ���� � � � � � �                 � � � � � � � �Ii�@
@   ��9����@� ����     ? H@    0? ���@`��         `����� � � � � �         4  ��0� � � �(��@      ��    `B ���    @� �AÁ�����&� �      �@    ����p� ��@��      3"@ ���e� � � ��`�+{foIo-�,n%�|��� � � R � @   #�/���em��+�֥� P J � % � ) P  0     �   � ��0� �@������� 8 p@ P@@p@`` ? ? @ `  @ @@"   P@��`����&� �0�@���  @ 
  Hj ��� �@�� �;��e � {��@�H���� � � � � � _ � e � {��@�H���� � � � � � _ �   @ �     � A < �@���������A�4���k#Ճ��GnC샯 ���x�����p��������+9��-�E��>�}> �     � +�QPџ�>�?����������`�� � ��`ବ�������   S    �� �	���yp���?�?��O���?�~�^�X�4�{�� � � ���	w@bxbx��&p�0� � � ���@�p�p�4��^� � ��> ~ � � ������������$ÜK"�r�_ ��x|<�<�������O�@s`�h_0,	���i(����������W������ � �Md-����i(>�?�d��wW������<��E-���i(������W�����PGC��]��'_������x�����C�� 4���(��:;��    � � � � �$�-�l�Hj�k٫�8� �� ���� ��y�����¿��0�A��y���g�/_0�p��б�!DȀW���_F�N�߀�����xȰ�ba�yx�@�>����a�a�y	��>�Qn��F� �
�"��&������������7�
����?�<� �~~ ������S@I b9�
�g�? ��������g8 �D ��q D � �- ���m��������?�?D ��q D � �MA[��m�������������D ��w O��������m��������   S@A<Br�y��1��xg������Q��1��f�                                � ���J �y,�ߞ����ƽ������zg��� ���D� ����q�s�g��_C���h}rXs�w�=�s_����������������8�-�o��W~��� ���������/���?�	�&"��
�F����������������vc��먥�od߀��{��{;�W�c���h}`Zq�w�=�s_����������������8�-������8�0����/������/��?�	�&"��
�F����������������vc��먥�od߀��{��{;�W�c���h}`Zq�w�=�s_����������������8�-������8�0����/������/��?    ����@�@�`�`    ������������
         � �@��@@���    ������������                                    P0!`BA                      �                       � @�����p                                      B�$Fqb!"AC! f               9�t@���		              �@ � 0�,@���    �          �` 1 0              HL�d! 0�R�  @             
����$%e!                    � @� ���                                     !!3����            !       /	DFF��            @        ( `��               �       �%�%�%�%�%�%�%�%�%�%______________________�%�%�%�%�%�%�%�%�%�%______________________�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____________�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____________�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____________�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____________�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____L
	
	
KM
________�%�%�%�%�%�%�%�%�%�%�%�%____KK________�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%______�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%______�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%L
	
	
�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%______�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%______�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____L
�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%______K�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%______KK
�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____L
K__�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____K________________________K________________________KK
__�%�%�%�%�%�%�%�%�%�%____________K____�%�%�%�%�%�%�%�%�%�%____________J
KK
_____6748944440____________�%�%�%�%�%�%�%�%�%�%_044:;4444@____________�%�%�%�%�%�%�%�%�%�%_0898944440__________�%�%�%�%�%�%�%�%�%�%�%�%_@:;:;4444@__________�%�%�%�%�%�%�%�%�%�%�%�%_6�1�2�1�2�1�2�1�2�6�_`a______�%�%�%�%�%�%�%�%�%�%�%�%____________bc______�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%____________________�%�%�%�%�%�%�%�%�%�%�%�%____________________L
	
KM
____�%�%____�%�%�%�%�%�%�%�%�%�%�%�%�%�%KK____�%�%____�%�%�%�%�%�%�%�%�%�%�%�%�%�%	
KM
__�%�%____�%�%�%�%�%�%�%�%�%�%�%�%�%�%KK__�%�%____�%�%�%�%�%�%�%�%�%�%�%�%�%�%K__�%�%____�%�%�%�%�%�%�%�%�%�%�%�%�%�%K__�%�%____�%�%�%�%�%�%�%�%�%�%�%�%�%�%K__ %%%%____�%�%�%�%�%�%�%�%�%�%�%�%KK
__%%%%____�%�%�%�%�%�%�%�%�%�%�%�%K__________%	%
%%____�%�%�%�%�%�%�%�%�%�%�%�%KK
__________%%%%____�%�%�%�%�%�%�%�%�%�%�%�%__________________ %%%%�%�%�%�%�%�%�%�%�%�%__________________%%%%�%�%�%�%�%�%�%�%�%�%__________________%	%
%%�%�%�%�%�%�%�%�%�%�%__________________%%%%�%�%�%�%�%�%�%�%�%�%___61212126_________________________04444440_________________________@?989440____________�%�%�%�%�%�%�%�%�%�%__67E;:;44@____________�%�%�%�%�%�%�%�%�%�%                                                                                                                                < B<�f�f�f�f�<<� $|8<<<�<<�< B<�F�>~ �~~�< C<�f~�f�<<� >~,�L�~��~ �~�`�|�f�<<�< B<�`�|�f�f�<<�~ �~�f~<��< B<�f~<�f�f�<<�< B<�f�f>?�<<� 8p �@@�            � Z�(4>?>4��" u"�T\(>}*�DD�  � � � � � � ���������u�6�J�I�I�J�2�HU.�V�6�U�U�R�R�@�N�6�J�	�U�"�z� u�6�J��	�J�2�HU>�N�V�U�y��R�@}�z�F�u�	�J�2�Hu�6�N�u�I�J�2�H}�z�
�U�U�*�*�Hu�6�J�5�I�J�2�H�O�`�@�@�@ � � ��7�@�`��p � � ��7�@� �@�0 � � � �        �        �                   � �U��������� �U����;����u�u�_����3�����b�u�޾��3�����e�b?�_���/�����U�^>�_����#�����]�b?�_���3�����]�R?�_���!�����u�u�]���3�����m�R?�_�� �        �        �        �        �        �       U����������U���        �             � ���           � ���           � ���           � ���           � ���           � ���           � ���           � ���           � ��         � ���         � ?�?��         � ���         � ���         � ���         � ���         � ���         �  � ��         � ���         � �������       � �������       � �������       � �������       � �������       � �������       � �������       � �������       � ����     � �����     � ?�?�?�?��     � �����     � �����     � �����     � �����     � �����     �  � � � ��     � �����     � �����������   � �����������   � �����������   � �����������   � �����������   � �����������   � �����������   � �����������   � ������ � ������� � ?�?�?�?�?�?�� � ������� � ������� � ������� � ������� � ������� �  � � � � � �� � ������� � ��������������� ��������������� ��������������� ��������������� ��������������� ��������������� ��������������� ��������������� ���������������?�?�?�?�?�?�?�?����������������������������������������� � � � � � � � �                  �
;������P��hH�  �����������$                      ��������+g-C��R!�%��                           ��g�_\g�cf�� ?�-�<#`c����                        �`���!1C�`�`�    ����������E���������I�#��������{��� M �������縝�ŗ�%#�����������n� ����������kw��.������������c�=������������������������������������������������������������������������������������������������������������r!�6��������������O���������u$����������������    �� �� ��   �� ����� � � � �� �   �� �� � � �    �� � � � � � � !����0��__�� ����� � ��_�� � ���<� ����� ��� � �� � � � � ��}� ����x� ���@� � ��x� � � xG�������� ���� � ���� � ̃ɇۇ�Ƿ�����������������������������������������������������������N?�p"���i�x ? � ���? � ���P���� 3��s5�� � � �  � � � ��Ƥ̈xC�,��t�����? � � ��_ϯg�sf�m���CO??�����?��������������������������������������N��;Ж���2-�����@� � � � ��{5�U�J1�{e䵂�v� � � � � �� �2�g|L�G����@ � � � � �� � �������߿��������������������������������������������������������_����5_��r��-#���/����? � �����������?�?�������������������������k��K�������������������i���� ������n�� � � � � YF}��87 +�'� � >� � � � � ��?O/OW?��_�K���?��O��_�?�?�8���>�u������� �3����������������L�����������`����������������ɜ������������7������������������������������������������������������������������������������������������@��������������������
0@w������� �h�������������M�- �45�������2�����������������������������������������������������-'Q����������������<�5���Ւ� ��<]L� 7�� � � � � � � �7�1YԾ@�( �`� � � � � � � � ���`��`q?g�*�� � ? � � � � � d�3���������)(�?��7����(���?����[ǧo0��������?�?�����������������������������������9����8��   �� ������ � � �� � v���> � ``����� �� �`��� ��	v����-    �� �� � � ��� x�����$ �  �� �� � � � � �� � ������ � || ���_�?� � �|�� B� �    �� � � � � � � �� � _���3s�0 GG� � � � � � �G�� ���?���   �� ���� � � � �� �         







     'O?\?Y>    �  ����� �� �  ����� ��     Z<Z<Z<Z<Z<Z<Z<Z<                                                                 � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U              �                  �<�~=�b�j�`~=�j�b~=<A � � U U �|��}�b�j�j�b�}�b�j�e` � � U U �~��~�a�j�b�}�a�j�`�~~ � � U U �<�~=�b�j�b�~�b�j�j�bb � � U U �|��}�b�j�b�}�b�j�j�bb � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U �<�~=�f�f�foM<�~��~~ � � U U ��<Y|9<�<�<Y<Y<�<�~=<A � � U U � � U U��~�~�~~�IU � � U U � � U U � � U U � � U U � � U U �<�~=�f�f�foM<�~��~~ � � U U ��<Y|9<�<�<Y<Y<�<�~=<A � � U U �b��b�b�j�j�b�b~�~�<YE � � U U ��<Y<Y�<�<Y<Y<�<�<YE � � U U ��<Y<Y<�<�<Y<Y<�<�<YE � � U U ��<Y<Y<�<�<Y<Y<�<�<YE � � U U � � U U�>�"�b�j�f::E � � U U � � U U>���F�V�F�F>�F~�<A U � � U U<�~��b�~�`�b~=<A � � U U � � U U��~�~�~~�IU � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U�<�<Y~�~~�<YE � � U U �b��b�f�l�z�u�y�l�f�bb � � U U ��<Y<Y�<�<Y<Y<�<�<YE � � U U � � U U|��|�b�b�j�j�bb � � U U � � U U>���F�V�F�F>�F~�<A U ��VV?���F�V�F�F>>A � � U U � � U U<�~��b�b�j�b~=<A � � U U � � U U|��|�V�V�V�V�VV � � U U � � U U � � U U � � U U � � U U � � U U<�~��b�b�j�b~=<A � � U U ��M<Y~��~~<Y<�<�<YE � � U U � � U U � � U U � � U U � � U U �|��}�b�j�j�b�}�b�j�e` � � U U � � U U�>�"�b�j�f::E � � U U � � U U|��|�b�b�j�j�bb � � U U ��VV?���F�V�F�F>>A � � U U � � U U<�~��b�b�j�b~=<A � � U U � � U Ul��l�q�e�j�j�e` � � U U � � U U�>�"�b�j�f::E � � U U ��VV?���F�V�F�F>>A � � U U � � U U<�~��b�b�j�b~=<A � � U U � � U Ul��l�q�e�j�j�e` � � U U � � U U�>�"�b�j�f::E � � U U � � U U � � U U`��j�e` � � U U �b��b�b�j�j�b�b�j�b~=<A � � U U � � U U|��|�b�b�j�j�bb � � U U ��VV?���F�V�F�F>>A � � U U � � U U<�~��b�~�`�b~=<A � � U U � � U Ul��l�q�e�j�j�e` � � U U � � U U>���F�V�F�F>�F~�<A U � � U Ul��l�q�e�j�j�e` � � U U � � U U<�~��b�b�j�b~=<A � � U U � � U UF��F�V�V�F�F::E � � U U � � U U|��|�b�b�j�j�bb � � U U ��VV?���F�V�F�F>>A � � U U � � U U � � U U � � U U � � U U �|��}�b�j�j�b�}�b�j�e` � � U U � � U U�>�"�b�j�f::E � � U U ��<Y<Y<�<�<Y<Y<�<�<YE � � U U � � U U�>�"�b�j�f::E � � U U � � U U>���a�e�j�`>>A � � U U � � U U<�~��b�~�`�b~=<A � � U U � � U U � � U U`��j�e` � � U U                                                                                                                                                                                                                                                                                                                                                                                                                                 � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U �<�~=�f�f�foM<�~��~~ � � U U �~��~�a�b�|�foo��f~=<A � � U U �<�~=�f�fo�Mo�f�f~=<A � � U U �<�~=�b�j�h�a�f�j�b>>A � � U U �|��}�b�j�j�b�}�b�j�e` � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U Ul
m
mJlJl
m
mJlJl
m
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
[
�
j
jJ�J�
j
jJ�J�
j
J
K
J
K
J
K
J
K
J
K
J
K
J
K
[

L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
O

J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
O
L
M
L
M
L
M
L
M
L
M
L
M
mJlJl
m
mJlJl
m
mJlJl
m
mJlJl
m
mJlJl
m
J
K
J
K
J
K
J
K
J
K
J
K
jJ�J�
j
jJ�J�
j
jJ�J�
j
jJ�J�
j
jJ�J�
j
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
L
M
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	J
K
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
�	�	L
M
_'p'u'v'u'v's'_'L
M
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	J
K
p'z'y'z'y'z'y's'J
K
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
�	�	�	�	�	�	�	�	J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
�	�	�	�	�	�	�	�	L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
_'p'u'v'u'v'J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
p'z'y'z'y'z'L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
�	�	�	�	�	�	�	�	u'v'u'v'u'v'J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
�	�	�	�	�	�	�	�	y'z'y'z'y'z'L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
_'p'u'v'u'v'u'v'J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
p'z'y'z'y'z'y'z'L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
�	�	�	�	L
M
L
M
u'v'u'v'u'v'u''J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
�	�	�	�	J
K
J
K
y'z'y'z'y'z''_'L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
_'p'u'v'u'v'u'v'L
M
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
p'z'y'z'y'z'y'z'J
K
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	L
M
L
M
u'v'u'v'u'v'u''L
M
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	J
K
J
K
y'z'y'z'y'z''_'J
K
L
[
 

 

 

 

 

 

Z
M
L
M
L
M
L
M
|'v'u'v'u''L
M
L
M
[














Z
J
K
J
K
J
K
_'|'}'~''_'J
K
J
K
mJlJ�J�J�
�
====�
j

0J 

 

L
M
mJlJl
m
mJlJl
m
mJlJjJ�J�J>�
�
>>>>�
z

3




J
K
jJ�J�
j
jJ�J�
j
jJ�JjJ�J�
�
�
�
====�
j
1
 � 


N
L
M
L
M
L
M
L
M
L
M
L
M
zJ�J�
�
�
�
>>>>�
z
 �


N
K
J
K
J
K
J
K
J
K
J
K
J
K
m�gJ�J�J�J�J�J�J�J�Jg
m�__
N
L
M
mJlJL
M
L
M
L
M
L
M
L
M
�m�uJtJuJtJuJtJuJtJm��__N
K
J
K
jJ�JJ
K
J
K
J
K
J
K
J
K
O

 

 

 


N
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
J
O






N
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
l
m
mJlJl
m
mJlJl
m
mJlJl
m
mJlJl
m
mJlJL
M
L
M
L
M
L
M
L
M
L
M
�
j
jJ�J�
j
jJ�J�
j
jJ�J�
j
jJ�J�
j
jJ�JJ
K
J
K
J
K
J
K
J
K
J
K
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
�	�	�	�	�	�	�	�	�	�	L
M
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	J
K
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	_'p'u'v's'_'L
M
O

__������������������L
M
p'z'y'z'y's'J
K
J
O
__������������������J
K
u'v'u'v'u'v'u'v's'_'L
M
������������������L
M
y'z'y'z'y'z'y'z'y's'J
K
������������������J
K
u'v'u'v'u'v'u'v'u'v'L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
y'z'y'z'y'z'y'z'y'z'J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
u'v'u'v'u'v'u'v'u''L
M
�	�	�	�	�	�	L
M
L
M
L
M
L
M
L
M
y'z'y'z'y'z'y'z''_'J
K
�	�	�	�	�	�	J
K
J
K
J
K
J
K
J
K
u''L
M
L
M
L
M
L
M
L
[
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
'_'J
K
J
K
J
K
J
K
[

J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
J
K
L
M
L
M
L
M
L
M
L
[
 

L
M
L
M
L
M
L
M
�	�	�	�	L
M
L
M
L
M
L
M
J
K
J
K
J
K
J
K
[



J
K
J
K
J
K
J
K
�	�	�	�	J
K
J
K
J
K
J
K
L
[
 � � � � � � � � � �L
M
L
[
Z
M
L
M
L
M
L
M
L
M
L
M
L
M
L
M
[

 �mJ�
�
�
�
�
�
m
 �J
K
[


Z
J
K
J
K
J
K
J
K
J
K
J
K
J
K
 

mJlJ�
�
�
�
�
�
l
m
L
[
 

 

L
M
L
M
�	�	�	�	�	�	�	�	�	�	

jJ�J�
�
�
�
�
�
�
j
[





J
K
J
K
�	�	�	�	�	�	�	�	�	�	 

zJ�J�
�
�
�
==�
j
 JJ 

 

L
M
L
M
L
M
L
M
L
M
L
M
L
M


lJ�J�
�
�
�
>>�
z
1� J



J
K
J
K
J
K
J
K
J
K
J
K
J
K
                                                                  %%%%%%%%%%%%%%%eeeeeeeeeeeeeee    %"!$!&!(!*!,!.!0!2!4!6!8!:!<!>!@!B!D!F!H!J!L!N!P!R!T!V!X!e    �#!%!'!)!+!-!/!1!3!5!7!9!;!=!?!A!C!E!G!I!K!M!O!Q!S!U!W!Y!�    ������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         !`  	     '                                             �� ( $$	$$$7                                                 �������'�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ?                           � � �                                                         � �                             ?                        � � � �                             ?                        � � � �                     � � � � � �                     � � � � � �                  � � ����  � ��  � � ����  � ��     0�?�?�<�<  �  � � ����  �  � � � � ��  �  � � ��� �  �  �<�<��?�?�  � � � ����0� �?����?�0�� �? ����  ��  � � ����  � �� ��������   ?                             � � �                                                         � �                           ?                             � � � �                        ?                             � � � �                        � � � � � �                     � � � � � �                     0 �0�0���0�0�00                  ??<�?�<<   � ������<��� 







                                                                                                                                                                                                                                                                                    <<bbbb``<<                bbbb<<              <<bbbbbb~~bb    bbbbbbbbbbbbbbbbbb          4444              ~~``````||``                ````~~                                              ||bbbbbbbb||                ``````              <<bbbbbbbbbb    bbbb<<                        bbrrrrzzjjnn    ~~ffffbb                                                                                                                                                                                                                                        bbbbbbjj~~~~                vvbbbb              <<bbbbbb~~bb    ~~bbbbbb                        ~~``````||``    ||bbbbbb||bb````~~          bbbbbb                                              0 0<     
                                       0 0<     
   @��:��ƭ���|� À���;;7�7�  � � @����@�@�`    � � � @ ` ` ǿ�;��·��� ' À���..-�0���������@�� �   � � � � � �                                                                                                                                                         bbbbvv~~jjjj                bbbbbb              <<bbbbbbbbbb    bbrrrrzzjjnnbbbb<<          ffffbb                                           ( -D<C(<     ?*                                       ( -D<C(<     ?*      9��C��w�C�d� �xCx{xwpsp||  �������`�� �   � � � � � �     4 � �@� �p�@�d|  � x@xxxpppp||                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    � @   � � �H�L     � � � �0�P�                                      3 O O$        � ��D<r��<����  �y��� �lx �`�� @ �@�     �������� @                                             �?�F����xa�� �������������                      <<bbbb``````                bbbb<<              <<bbbbbbbbbb    bbbbbbbbbbbbbbbb<<          bbbb<<              bbrrrrzzjjnn    ~~ffffbb                        ~~``````||``    ||bbbbbb||bb````~~          bbbbbb          ������� ��� � �� �� �    �����                                F#s3<   3    ��=� ��� _C䟌{9 � ��8  ��{�s{                                                                                                                                                                  �                                                               �                                                                       @ � �                                                           @ � �                                                                                                                    0 0                         ||bbbbbb||bb                bbbbbb                                                                                                                                                                                                                                                                                                                                                                                                      �                                                                                     bbbbbbbbbbbb    ~~``````||``4444          ````~~              ||bbbbbb||bb                bbbbbb                            � ��`@� Ѐh��d    � @� ���@��                                    7U^H        <? | � � bd��w� @   | ��g�`  �� �   �@��@��   ��  ����                                        >*=
            �|���~N2���< ��������r�                                    �                                                               �                                                                       @ � �                                                           @ � �                 $�����|��`� � ��p� `  �`                                    g'/	  ;   �����1�|��!� 8�������??��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 0 0                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                                                     $$HHllll                                        <<bbbbbb~~bb    ~~bbbbbb                        ~~    <<bbbbbb~~bb          bbbbbb              <<bbbb``````    bbffllxxppxxbbbb<<          llffbb              6666$$                                                        ||bbbbbb||bb    bbbbbbbbbbbbbbbb||          bbbb<<            ` 8@()

       (   	               ��                 �p�x�4�*C!
 �0�X�$�}>             ���@`           ��@@�  ) "!UCVA   ????  ��pp�(�d���.�   �������������    I6K7V/         	  P   �`z��l�x��z��@     � �   >  !	 	
   1       � �P� F�N  � � � � � � �  ya���Osc��sc  ~��������|  �8�������  ��~��������~� 'x0`5uA!  0 8 O J j ^ � (��XH�>������� X   � V V z                                 56� 	

+*�                              ����PP((
                                      �.@�6 x � � � G ���0H@�D�B� GIDND)&&   ????   R�F�Lpp��  ������������ �  �z?���v:4        � s ?   L�耘 X 0 � �   > | � � � � �    14t{X|~~~~||�  0px~ ~ |  � � `d�          � � �         8p0�@�@�0h����������������8���w"g20* 0   H H j ? *     ���輨T ��( p     V � | � �   /DP�B�!�,M >3 | �C�?�s >P(�� ^� C �   � �(�D��g � �      ~~����Oo:;    ~~����;;    >>��K�����Pp    >>��������pp   8 <.&&   ( $ " " "   
/^,�$��@   ) R � � <    !+_ _      ?4x}   � p�����0�@�   � ���(0�0��<  ) "!UCVA   ????  ��pp�(�d���.�   �������������                                 ��� �           ��� �                                    x �h%6�           �                                  � V "�T          �$$p�            	                      � ��            L�N
<$ld8800<<\|(800Hx$<

||00xx<<l|0076    	    !     �@�@�`d  8 �   8 < � � � � �   O/'     | ? ?       �Đ�p� � ` �    �<�|@� � � �    IDND)&&   ????   R�F�Lpp��  ������������ �                                                                               +6Qb���x�����pr � �> > ���p                � � �"#������pt ����܈$ ��� t   		      ����\������LH P� �             �>                  � ��`@x`.���      @�����p�:�j^<~{3/~~_;?? <<~��?0~��@                                j^<~{3/~~_;?? <<~��?0~��@                                                                                                   @@D        PPDD         @@D        PPDD        \T)  @H01@H
^))"&   @@D        PPDD            !  0  PP	L\

!!Pp$$  \T)  @H01@H
^))"&      !  0  PP	L\

!!Pp$$   @@D        PPDD      �pz     ?       W֯��������     :�������                                                                                                                                                                                                         @@D        PPDD        \T)  @H01@H
^))"&   @@D        PPDD         @@D        PPDD         @@D        PPDD         @@D        PPDD         @@D        PPDD        \T)  @H01@H
^))"&   @@D        PPDD        \T)  @H01@H
^))"&   @@D        PPDD            !  0  PP	L\

!!Pp$$                                  
,4<$0h 	 	  " B B �      0 	 
   $ ( H                                  &`��� .P     H v                                                                                                                                                                                                                                       @@D        PPDD         @@D        PPDD         @@D        PPDD         @@D        PPDD                            p8(X `�� � �    � � � ` @ @ � �   @` `          P � � `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          9G?�r�Y�mZ%_        $       � ��4�����b��`�      p      f0ad?�g�w�`�A�1 ?00xppxwxG � ������8� � � ���H��� �� < 3 �06����`��   � �0 ��`��E��`�8j�� � � `x 4��8 � � �`v��zo���@p  �� � ~>�� @                                 #g,s(             #g,s(             #g,s(             #g,s(                                                                                                                                            @%:::* .  ?       v�LԨ�x�0�� � � `����� �    �p� M^?- {~ ys? ? 11>>  P�P�p��@�`��    � � � @����    ��|��b��   �8�8` �   h���H��@��� �@� � � �00p �  ��  h���4��� ��    � � � �  xx                                     #g,s(             #g,s(             #g,s(             #g,s(                                                                                                                                            M���W������� L��� ���� �M���W������� L��� ���� �M���W������� L��� ���� �M���W������� L��� ���� �                                                                                                                                >5{:Fo0�k�W�N            `X|�ڴ~TnԲL|���     �        \=0(#j;U5K)])    
 �x���Vܪ�Ҕ��� �`    P h@h( �
;������P��hH�  �����������$ sP���
  #�gW�G�(�$�                                                                M���W������� L��� ���� �M���W������� L��� ���� �M���W������� L��� ���� �M���W������� L��� ���� �                                                                                                                                R<W8/10      F�f � v�������� � � �,�,��  �ge6�Ed?%?, A /  �Цl_�&������$�(  � �`�`� � ���������+g-C��R!�%�� !1o_���������/J��  ( �(���8                                                                   ��� 	[  0       @ @ U�  AF	                                 �  �"                       ((      �QT  D  �  &    �0�0@c � &@7  Ft  Ft  �9<�4�4jtjt    `@`@   @2    ���  ���   F�       �    � �X� =	�
  \�� \��     iv������� ��UUUU��L UUUU�U��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� �L�~ /�mJJJJJi��'''�  ��_D~�Y�~    &   �8�n�n+m��`i�e�e  ~'c�  '� ̰r�UUUUUUUUUUUU�ܤUUUUUUUUU�!WUUUUU UUUUUUUUUU�4�>� UUUU� �   UU�      �  "                ! �  UUUU�1����	� �    � � A) �    �  >   �UUUUU  0%�����    � B  �� e            +'���##���+ !�)�  }�#  !���~� �   � �Z�>�c����ӳ�����£�C�%K��������k�*���k� �U�h�R�$             IHUU   UUUUUUUUUUUU      UUUUUUUUUUUUUUUUUUUUUUUUUU     
     O   �                   ��   �         D�  �� �  ��             @ �                 [Gs�aW3]�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU 0%������ � B��� Bc�$ B'��   B��  ��" !���~  
         UUUUUUUUUUUU   p � � � ��������UUUUUUUUUUUU    UUUUUUUUUUUUUUUUUUUUUUUUUU  x �UUUUUUU  P%���   ���_ _�/P_ _�/0� B %���_ _�/0$ B5�� Bc�$ BԢQ �  �����~   ��   �	
  "Q� "0� 	      �   ,�    PR�s     ,|          ��e	���  j/=�0N
��Hm,
��e�%�O�gF��H�!m,��eO��hF� H�!m,��eO��L
�� @�-k%J!��O1�4��gF��` �e	�=�5�5K/=�0M�gF��` N-��B f�$�$` ) 1e5�=�$�c)%J)k-�1�5�9�=B1FRJsN�R�V�Z�^UU���<1!�-�B�df�Ip^0s�|�UU�t��U.W�6�W�8]]_vS`9�{UU�� z5]>�::WCr�-�6�[8U�z�UU�w�f-�-J?�G��j ��R�1�QR  ,��S��f{�z�Uv�~/~�	��5�� ��5�R�yZr�~]5�.^7�_��� ��5�R�yZr�~]5�.^7�_����3��h<��j<��l<��n<�� 2��D1��F1���3���#�� "�M
3 �5 �7�@3�@s�P��P�H�8���8�� 2�� 2�� 2��>��>��>��>�� 2��@:��Bz�� 2�� 2��"��"��"��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UU��UUX��3��h0��j0��l0��n0�� 2�c�3�s�#�y ",Y�p<Y�p,i�p<i�p8h 2@p
B0 2�� 1�� 1��&1��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ��UQ                                                                 	
����������	M(              (              (                                                                    UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� ����
��! ���0)?�:ȹ ��Z�:��! ��z� ��:�� �`�� �  �$  �rUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���������������������������������������������������������������T	*:	)5����������������������������������������������������  @`�����'�N�' O ��g� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �`"�"�"�" ��" � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �`````` ` ```````@` `````@````` ``` ```````@````` � � � � � � � � � � � � � � � �`p`p`p p p`p`p`p@p p`p`p@p`p`p p`p p`p`p`p@p`p`p � � � � � � � �� ��� �� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �@���  `� 	���������������������������`�������`���`���������@����� � � � � � � � �`	��	� 	@	�	�	 
����	 
����������������������`�������`���`���������@����� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �                                                                                               * * ( ( ( % % % % # # # # ! ! ! !                                                                  �@�[�o�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  � � � �  r h _ W R L H C ? ; 9 6 3 1 / - + ) ( ' & % $ " !                                                                      
 
 
 
 
 
 
 
 
 
 
 	 	 	 	 	 	 	 	 	 	 	 	 	 	 	     �������������	#'*.269=AEHLPTW[_cfjnruy}���������������������������������� "&)-158<@DGKOSVZ^beimqtx|������������ �~H � � � � � � � � � ~ w r l g c ^ Z W S Q N L J H E C A ? < : : 8 6 6 3 3 1 1 / / - - - * * ( ( ( & & & & $ $ $ $ ! ! ! !                                                                UU �F�`�s�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  � � � � { o e \ U O J F A = 9 7 4 2 0 - + * ( ' & % $ # !                                                              
 
 
 
 
 
 
 
 
 	 	 	 	 	 	 	 	 	 	 	                    �������������!%),048;?CGJNRVY]aehlptw{����������������������������������
 $(+/37:>BFIMQUX\`dgkosvz~������������  1        2�      ��  � l $       � c T    P} �|�y�X�    v���r    �~�~�   jՙ�    � l $              g#V����������|G}J~M�s����                                 � H �8  ,      � � �8       R�F�Lpp��  ������������ �    ) "!UCVA   ????  ��pp�(�d���.�   �������������IDND)&&   ????   R�F�Lpp��  ������������ �      ����       �RUY���Ѐ��       ����    ������������������������������������������������������������������������������������������������������������������������������������������������- - - - - - - -                                                                                 ������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                ��������������������������������������������������������������������������������������������������������������������������������Q�  I�       g                                                                                                                                                                                                                                             )  � �    � ��X�                                     �M�]�w����ݑ'���׻��e��y�d�      �:�r�J�5��[�                                                                                                �     �M �    �`��� ���@���@�`�`�� �`�pUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��;��w�ݑ���]�`��Պ�MgY��Պ����׻��MQeܠ����y�R�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU        5O             �               �            �   �           ��         �  �          P��P�        �    �            " " " "     " * "                                                                      (4h���    2 B �     0 `   	  $ H � ``@�            �   �               0     	  $ H p @���              @ �                 (8        4 �   $<��� ����   1 �     @ �                        	     (@� �      1 �  ` �   ����             ` �             
,4<$0h 	 	  " B B �                       p8(X `�� � �    � � � ` @ @ � �      0 	 
   $ ( H   @` `          P � � `                  " " " " >6   A I "          ��      �  �         �0���0        �    �        �  _   +      �  _   +   � ������   � � � � � � � w>*>k6w A   A c c w k   ] U\" ] U  T    6       > q G � �       > q G � �         �  f M         �  f M � � D "         � � D "         H D             H D                                     � @ � �   P �  � @ � �   P �                      0 h � �   p � 0 h � �   p �                                     ~ � �         ~ � �    � �  � � �    � �  � � � t �     �     @ t �     �     @    1 " @  �    1 " @  � � } �   "     � } �   "     � � � c �      � � � c �        �   �           �   �                 p �          p �     � �  ? �     � �  ? �   � � � � � � �  � � � � � � � �     �     �   �     �     �                                p            p           �  �  0       �  �  0         �   �           �   �              
             �@��` `      �     �     
                        @�� ```        �  � � `           	                    ��0�pX8,      � 0  � B  <,0          4 @ @ <         <8          "   8         < d�� �{���$  8 p F b  b B �B� �&{���|<$ f @ & r $      6 n �8�V ~v0   8 @ ( 8 (  ~V.h^~^x8( (  0         < t�
� ;��@{  8 t f f &  
 ; ^ �$�@�"�P?@?  8 P   \ .     < t�
� � _�{  8 t f f &  
 �"�@�
�|<  D & t (        + � �D    
  > V " ���(� c   d o W        z�D�*� � \�� �  : T ` `   | j � �#�@�
�|<  D & t (     < t�
� � �@�]�  8 t f `   | * � ��"��
�|<f b D & t (     ��D�
� � � z  : t f F   
 ' >> 0,>            < t�
� � �@��  8 t f f & < ( �"��"��
�>A> D b D & t (     < t�
� � ]�� �T  8 t f f " f * �#;B�@�
�>@<    & t (             8Z � �           < ^ f ��� � �
�<C<d b F f t 8               .|            8 v 6 >".>>                     < @�#�          < \ b � 4~ �"�Po'   0 \ .             < D�*�           8 T f � "} �D�#�?@>    " \ 8               *h             �� ��&z�w  h L n X               ~��@�"�          > \ ` ������$|"t n  B |              > 
A� �           < ^ ` �_����$� ?@> t . b d Z <             ~��@� �          > ^ d � }?,2, <   
                 < Xu��           <  f �@^�� �� [�~<& 8 f d ^ <             8~;��          8 v f � �@w�?��`�|<f >    ,      n � ��D� P<    f d " f ,    0l 4 (0,     8        j <�{ 3~ _�?@   f   0 :    v� |� W"  , F   f ,    &`��� .P     H v    :D�� >�� l#<  z ` t  f    <*`�@�_��Z 8     t & d <   v��Cz 0(<    v $        x"� nJ�� @<    f 4 b F <   < v��D;h= ^<  , d "   ,   �0 0�� �        � �                                        ���`p�0�          � � �                     ��0`p�� �      � � �                00                 ���08���        � � � � 00                 ���08�� �    � � � �            00/`/`              ���08����      � � � � � /`/`00              ����08�� �  � � � � �                                        x � � ��� ? H0�x���8               �         �    � � � �  @?����p    � � ���@� �	 ���� � �  	        +         $    @ � ? �@  ��<��  �������  � ������           � 
 �          �
 �(�� �� �D� � �(�� � � � � �8�| � � ��� | |D|88�|�|�|�| |D8D88   ��$<��((    � <  � ( !!��!! ! � ! ��@�(� �B�HH �@� � � � �@H pp������uw p��� � w�@@         @     <<``����������B~< ` � � �0�� ~�b~<<        ~ <B             ��  00      �   0                 ��           �  ,<�� �    ! <@� � ���p@0?��p(?�|t>A� != � � � �� ��� � ������p�                       ���            � �                                     � @ `   0 2Hy���  @`    "i�         	 A ��� � ��   @ �h`� � ��  �@��``� �"> �@6   x���� �                            ,=��*���@� � � =�@�A��x��_��  ��@@@@00�   � @ @ 0     ����     !� �  � � � � � �     � � � � � �       � � �  � #    � � �  � #  �   @           �   @                 	        	  � � � � � � � � � � � � � � � �             �             � #  �   �     #  �   �                       � � � � ���@�?����?�?`                   q��0�    � 8�� �c ?  � #@'   @���������p��8�� � � � � � � �    88(((   88((((((((4 4 ��(((((  �     088 0   08 8 0((     ?�|g??         ? |�?@ ?    ����   ����   ( ( ||((((( 8 8|�800  "!	          � @����       ��@@��P�h3
 )

 �BF,(0       B�z$0 0            (8           8 /        ��     ���   lD(((( (T|( |D8(((T(T| (| |D| 8       | | | 8        88TDlD8XXh0(08DD8D8(hl0L0LHpHp0(0       pp00                
	                ��  � $�        �  � ��$#                     P� ��@    ��    � �@� � ��                       �
��         ����('PO��           @?�          � � ��@@ ��``   � � � � �@`     ``XX0 &(	  ` X        d�`� �   x � � �	&(0 XX``       X `    ���`d   � � �x      ��      >�|   @@$   $ ��@   > < < |� ��  $   $   ���  f ~ < < ~ f�    UI   H     A>  H� @    *"  HH��@@    " H �@@   """"      " "                                                                   �              @ �                          �                � @                             ?      � �``�`� �     � � � � � �
        ? ? ?       �� � ��        � � � � � �          `   ?     �  � �  �,�,�T�"� � � � � � � � �@?@?@?$*      � � �   ?   ������pp    � � � � � � � p   	     b "@      c � �  0 (        0 x � <  '   @`        � � g 3 < > >    �     p    8 � � �  x � p           @ @   <      @ � �               0 8     @                   @       1 0                               p `                                       � @�             � �                           @��              � �                                                  � @�           � � �                          @��              � � �                  
	                 ��  �P�        �  ���
	                 P��  ��        �� ��               	
	             ��``�P�(�      � `����
		             (�P��``��      ���`��           ('('           ��00�(���    � 0�����('('           ��(��00��    ����0��       ,#('POPO     @?@?  ��00�4��
�
�  � 0������POPO(',#  @?@?     
�
��4��00��  �����0��                                   xx������??0xx������'?     ��        ���������xx  ?�����p�  �����������������@� �	      -)        &/    �?�����?  ���#?���  ��������������  ������������        ��*
��        �� *(�� ((���������������� �� �D�8�|�������||||||88  |�|�|���||8|||88              ��$<��((      ##��##  @ ��������@   ��`�(� �b���HH� zx||vv� ����������                @@            p@B@\\�<<<``����������B          b~~~                            ��  00                         ��%(P  ��� ;?6>l|��0���??O__#��sKq��p=?*?����������������������������r��                       ��              ���                                 ��@@@@  002211yy �@@ `   02Xy��     A  			CC  �@�  � �@���������������`�����  M�*>��    x���                    EՕ??������.?��k���P���_�                ��  ��@@@@00   -00    3?����������������    ������������      ��������##  ��������##��  @@          ��  @@          				��������������������������������          ��          ��##����    ##����                     ����������???����?���_             ������ q���0���aa  �Bc8?��        ������@���������p��8�   8<040$0$0$  <<<<<0$0$0$ 4 4<<<<<<<<<��   000000  (888(8(8(8    c�X ?         ?��g??       ��� �    �������  0000 ((� (8(8(8(8888888��  ,.
   882>1?      � ���`@@(      ��@�������%	   ;?,�8B4       ��~~,<(800            (          /? ??        ����     �����( l((  T |(((88||||8888||T|T|TT||8888      (| |D| 8       D (( ( H$HXT||||||88xx||l|l|484808      L|L|8(8       P�B���@�(� ~  ������������~~  qBq�1��  ?  1�1�q�q��� ???  !YH�D�  �  PP��������   � � ��� �  ������N�����  @3[0@(M9@-B8� !�!�1�0�(����E�ŉG @���`�E}�������� �?���D D D DHX �  D�D�D�D�L�P���  �D�D�@�C�"`1 �  F�F�B�B�c����  1@qFp0F " �� pc�#�"�"�����pp � � � � � � � ����������LLMO]�� �  NNNN�����  
�
���L�D� �  ��������������  �� c`�p�  �  a�a�������`���   "! 1�� �  ������������  �O�O�F�F�GF �  F�F�O�O�����   0 80  �  ��������  <Bb��f���fb�<B~ � � � � � � ~ "<DqI:'G��3��> | y ?  � � � ]c���4�b�@�m�;?� � � � � � � � ;J��!�q�s��>A]b{ � � � � �   ���|�/�f���� � � � � � � � =C&Y��������g��%  � � � � � � ?@��������`��|� � � � � � � � "<DqI:'G��3��> | y ?  � � � \b���4�b�@�m�34�~ � � � � � � � @>A������p�p��   � � � � � � ��~�,(XhxH0@0@� � < 8 x x p p *:I)!"@p`PqQ; { ; 3 3 p p q �(��}U���8â ��E� � } � � � � � ��m�E�KG����<"� � � � � � � > 0 0             0 0                                                                 >"fT2P ��E�A  > v r � � � �   ��g�g�~��D�L�  � � � � � � �   AY� ��@�@�ez   � � � � � ~   | �c�ŁG�J�  | � � � � � �   ���`�|��@�@�  � � � � � � �   ���`�~��@�@�@  � � � � � � �   A_>`� ��I�d~    � � � � ~   c!�B�|��B�B�B  c � � � � � �   " 8D  >      |    �J�J|      � � |   ¡�6�t� ��J�C  � � � � � � �   @�`�@�@� ��@�  � � � � � � �   F�G�+նm�Y�A  F � � � � � �   ��r�z��V�J�J  � � � � � � �   Zf�GŃ�Fj�4L  ~ � � � � � |   ��åg�k�z��@�@  � � � � � � �   < Z<c���D�Ft
  < ~ � � � � ~   ��åc�i���B�B  � � � � � � �   _a@#` zF�A��   c ` ~  � �   ~�sk8(8(8    � { 8 8 8 0 0   c�c�B�B��B�J|  � � � � � � |   ƅ�l*nthP(  � � n n | x 8   �C�G�E�d�V��J  � � � � � � �   A"cU*<$hTĪ�  c w > < | � �   A""DvZ$(Hx0P  c f ~ < 8 x p    0@ �       0 ` �               @               @             p   `          p   ` *:I)!"@p`PqQ; { ; 3 3 p p q �(��}U���8â ��E� � } � � � � � ��m�E�KG����<"� � � � � � � > x � � � ?�  0 x �                            �                   � � � � x   ?  � � p     � � � ��@� � �                   -                  ���  � ��             �������    � � � � �            � * �(         �     ��(�� �� �D� �             8 | � � � |�| | 8D 8| | | | | 8 8       �$  � (                 #�#                  @Ġ`�(� �b@� H                ��z�|�v���                      @                     < ` � �p�B�\���                bB~                             �   0                              �                 %;(6Pl ��0��                �p?@Op_�p#<(         � � � � �� ��� � � � � � p                              � �                                                      � @ @   0 2 1Hy�  @             AC             �  @@ ������`��  � �           �"     @        �x�                                           .E��j?��@� �          � _  �   � @ @ 0                    -30� �                � � � � � �     � � � � � �       � � �  � #    � � �  � #  �   @           �   @                 	        	  � � � � � � � � � � � � � � � �             �             � #  �   �     #  �   �                              � � � � � �?@?    ? ?                             �q��0          �   �a      @          �@ � � � ��p��8                     8 0000         000  ((�          (00(0 0                    c'            � @ ?       ����            �     0 0 0 0  0��     ( (    
                     ���@��@�@�             (    !         ,n8<         � B $               / (8                      ���        �     (8llT(88T||T(T   (           T(| 8D8                        D|(lT  0$4$Td   ( ( H H H  4D4D0                     < d�� �{���$  8 p F b  b B �B� �&{���|<$ f @ & r $      6 n �8�V ~v0   8 @ ( 8 (  ~V.h^~^x8( (  0         < t�
� ;��@{  8 t f f &  
 ; ^ �$�@�"�P?@?  8 P   \ .     < t�
� � _�{  8 t f f &  
 �"�@�
�|<  D & t (        + � �D    
  > V " ���(� c   d o W        z�D�*� � \�� �  : T ` `   | j � �#�@�
�|<  D & t (     < t�
� � �@�]�  8 t f `   | * � ��"��
�|<f b D & t (     ��D�
� � � z  : t f F   
 ' >> 0,>            < t�
� � �@��  8 t f f & < ( �"��"��
�>A> D b D & t (     < t�
� � ]�� �T  8 t f f " f * �#;B�@�
�>@<    & t (             8Z � �           < ^ f ��� � �
�<C<d b F f t 8               .|            8 v 6 >".>>                     < @�#�          < \ b � 4~ �"�Po'   0 \ .             < D�*�           8 T f � "} �D�#�?@>    " \ 8               *h             �� ��&z�w  h L n X               ~��@�"�          > \ ` ������$|"t n  B |              > 
A� �           < ^ ` �_����$� ?@> t . b d Z <             ~��@� �          > ^ d � }?,2, <   
                 < Xu��           <  f �@^�� �� [�~<& 8 f d ^ <             8~;��          8 v f � �@w�?��`�|<f >    ,      n � ��D� P<    f d " f ,    0l 4 (0,     8        j <�{ 3~ _�?@   f   0 :    v� |� W"  , F   f ,    &`��� .P     H v    :D�� >�� l#<  z ` t  f    <*`�@�_��Z 8     t & d <   v��Cz 0(<    v $        x"� nJ�� @<    f 4 b F <   < v��D;h= ^<  , d "   ,   k-�1�5�9�9�=BB1FRJRJsN�R�V�V�Z     !!!!"BBBCCcccdd������������ � � �~x��   ͍~x��       �    "�,O�~�d�   7              5   ��[ ț ���(�) �* ���+�+ �, �-��~�u�   ��~��    & 8 J \ n n n � �       

  �
  ��  ����  ����  ��  "9HW%RUN"9QbP)H|rX4Pa��n"2N[s���F[o|���P@��D� Bf�@@� D�Af�@H 1@HV  "& H !H V )& PP	LT

  P`$$ P 	 T
  !`$    P@          @ D         | �?|          ?�        � ��
����        ���� �      ""  666"*" """6                                t �0�� �        |0���`!P�|��       0a��< �      @ �              � �                                             ( p �`@`�      8 P`�@��  	  �@���� �       �`�@�@ � �                              j�0Xp(��  v0�p���0                      "D� ��`�6l ��0� `����           � �@ �                    � @ �� �`� ���`@ � ��@�`� � � @�   }�?}        ~?�~      � /��/��     ���� �  ��O tP_�π@ ���@ ��_��x�O ��@  � ������        ��~��~ �              `� � �`� ���@ � � � � � �`�@ � �                          � ` X����|       � ��8�|��0W=i�8�x0�i>w8�x�                  ��X�` �         ��8 � �         �  Y     , �  Y     ,     � � � | � ^     � � � | � ^ . � U U  U  
 . � U U  U  
                          �  `   A   �  `   A  � � �  �  �  � � �  �  �      � � � � & �     � � � � & � 
           
           0   `@ @�� ���  @ @ �@�@�@ ��� �`@ @0   �@�@�@@ @               
                        @��            � � ?;Zo��Uo=
8/nO��MO05
  ���^�����P\���� ^���P� \�� :4/Po��Uo=
 0pO��MO05
 P��\�����P\��� \����P� \��   0��Po=
  -`�@O05
   P���P\��  � �P� � \��    	  	            2P � � P 2  < p � � p<                      ��     � �  � �     ��        $  B B$f        < f f$B $ B f  � �B� �  < f f � �B�B�           $ B             < ff  � � �B�B� � � f � � �B�B�B�B�                                                                RPPRPPRPPRPPP  PP  PP  PP  PRPPRPPRPPRPPP  PP  PP  PP  P <b �D�B����@�< B<�~�f�f�f�f�f$�B� ل�b��>�f�f�f�f�~�< >  6n �"�(V nF &F8�x�8F8F8F8 n(FPF V f F~>F8F8F8F8F8F8~ >  <
r� �Ļ �y< B<�~�f�f�fy; ^� ��"�@ ?#F8�p�`�~�~ ?  <
r� �D���y< B<�~�f�f�fq {� �$��>y�f�f�~�< >   
1% R�� 	!A>�v�f �"�U� �ey  �f���y	  ~�� �@����"�~ �~�~�`�`�`�|�~ � {E� ���>�y�f�f�~�< >  <
r� �@� ��< B<�~�f�`�`�|�~@� �D���$��>�f�f�f�f�~�< > ��(�� �D� �y� �~�~�f�f�y' . >6. . > #&&&&&>   <
rD� �D� ��#�< B<�~�f�f�f�<�<@� �ـ�d��A >�f�f�f�f�~�< >  <
rD� �D�����< B<�~�f�f�f�f�~� {Dy �d��@~ <�>yy�f�~�<~ <         <$ZH� �        < B<�~�f!�@�D� �D��C>�f�f�f�f�~�< >          &~         &F8v6&&2.& . > f&&&&&>           <hVE� �        < B<�~�f � {
& ~�*�?�s&N0�~�~ ?          <`ZD� �        < B<�~�f�,1} ��3�@ >�1y�f�~�< >          0.TB         "B<`�� �@���w �l�L�~�~�s          ���@�!�        � �~�~�`@����$��">�|�~��F�~�< >          >uK� �        > C<�~�`P����!�@�$�@ >�|�~�f�f�~�< >         ��(��E�        � �~�~�f �y ;'*&, < �q#'&$<           <&Z�� �        < B<�~�f���"��D���>�f�<�f�f�~�< >         < zĳ#�        < B<�~�f �2������$�>�f�~�>��~�< >  <N �� �B�`N << B<�f�f�f�fB<<   ,l4$ ,,  $D8$$$$  <Jý{# ~��@< B<�fy#N0�~  <f� w}&�(G">< B<�Fcy�fC<>  2*`~H���P~ "r�L�~�~ D~h� ��� {$�O>~ �~�`�|y�fC<>  ,TJ �D���D�$Z<,B<�`�|�f�fB<< ~T��z ,$ < ~ �~�fr$$$  <ZB�$"�D�hV << B<�f ~�f�fB<<  <f%� �DS=!O>< B<�f�fA>9C<> UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�� 2DE ��$T�PP��EQ���  \T)  @H01@H
^))"&      !  0  PP	L\

!!Pp$$   @@D        PPDD         |G�|       ��       �0/��0/ �      ���������        **6>6>*>6*  6>">*>6>                            t@�@P��      ||����`�./Nh��� �      1?q��|���      �@ �            ����                                          ( P ��P��    88pp���`� ���� @ � �      `�@�������                             bX��(����~~����8�0�                      
*8TP� ��6>l|����`��� @ �          `�����                   ��@ @������@`� ������`�`� ����   |G�|       ��      ������� �  ��?��?��� @�O�s�s O�@ @����������������   �@>��@> �      ���������            ���������� @�@ �`� � �`�`�������                      ��`��HD8�      ����x�����\�(A< a\�4���??����                HD���` �        ��x�����        ��YY,,��YY,,    ������||��^^    ������||��^^..��UUUUUU

..��UUUUUU

                ��``AA��``AA��������������������    ������&&��    ������&&��

      

       0   `@ @�� @000`` `��@����� @��  `@ 0  @���@�`` `000                                     ��(�            @���7j.�5T]*:(*8?0?����u?
����*�{s]��PP�������������o?�?T]*:(*??p����u?
��,�����]��PPP������������  
(O/pp/?(*  ??p��p?
  ��T����PP  P���������        1 P@�@� P1>?pp����pp>?          s� �     �s�����    ����       $fBfBBB      <<ffffff $$B fÁÁ����<<ffff�����Á�           $$B          <<ff fÁÁÁ��������ff���������ÁÁ�                                                                 PR PR PR PRPRPRPRPRPRPRPRPR PR PR PR PRPRPRPRPRPRPRPRPR<<dx��߽�{���� <>~~�f�f���f�f�۽����{?����||<<f�f�f���~�<�>6>n~����V~~nvN >8~x�:�8~8~8~~nVn.^v~f^fxx888~8~x~8~8~8~~><<tx����;߿{} <>~~�f���f�;?^~��޾��ݯ?????8~t�`�~�~�@ ?<<tx������_?{} <>~~�f�f���{��������||<<f�f�~�<�>���� ??>v�f��������f���&�g  zz��������\<����~~�~�`�`���|�~���{��������||<<�g�f�~�<�><<tx������߿��]+ <>~~�f�`�`�}���������?����||<<f�f�f���~�<�>׻��������z|��~�~�f�f��'?>.>>08,<>.?>>>>> > <<tx������߿���� <>~~�f�f�f�=�?�������?����>>>>f�f�f���~�<�A ><<tx������];���� <>~~�f�f���f�~���{;=������>><<?�Ff�~�<�@~ <        88Z~����        <<~~�f�������������<<<<g�f�f�f�~�<�C>        .6||         >:~v~6> .6>.>>~>>>:>>> >         <<>����         <|~�f���{4,~~��կoo''�>0~~�~�?        <<:����         <|~~�f���}߻����??>>�.?f��?�@ >        *        <>|~�������z~wl�L�~�~���         ~~������        ��~�~�a�����������|||�~���F�~�<�">        >>
>����         >}~�`���_/��������??>>|���f�g�~�<�@ >        ~~׿�ߺ�        ��~�~�g���}{?;,4,<<<�??:>< <         <<X|u��         <>~��f���^z������[~~<<f���f�f�~���>        88~z;w��        <<~��g���Ϳw]?;���||<<f�~�����~�<�>n^����߻��.<< <<~f�g�f�f�|~ <l|4<(0,< 8<8|<<8<< j^<~{3/~~_;?? <<~��?0~��@vn��w|~��Wo <<~F�f�<">������.. >>l~L�~��P~::����>v{��l\<<D~~�`���f�?><,*ܼ��_?��Z~88<|~`�|���f�<~<vv����z~(0<<~~�g�~8<<< x\��n4����><< <>~f�~~f�f�|~ <<<vn��߻;=?^n<< <<~g�f�~?=>UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUF  |�s    |�s     ,|          ���%�B� �_~e�<*�%O���6x**�%O��O��3'�&�&*�f��\G�:X.�-n!��.&�R��&*� ��\G�:X.�-n!��.&�R�2*�)N! ��Z[�J�F:�-)�f�i\=R'�&�&*�F�����[ko�4_~e�<��&�&*�f����[���.����&���@�� V`b�j��IUU�w�f-�-J?�G��j ��R�1�QR  ,��S��f{�z�Uv�~/~�	��5�� ��5�R�yZr�~]5�.^7�_��� ��5�R�yZr�~]5�.^7�_�0�� )��  ����  

�� ) ����;i h(+`�0� �H�H�h�  _��� � �  �  �H ְh x֫(+`�0H;8� [�� �H�H�h�  _���� �� �� )� �� )� �J���e��� �  �����������<� 鬤�  � ��� 8�




�� � �	F� �F�  )� 

�e�� �� ;i	 (+`�0;8� [� ��H�� � �� _���� ) ��  )� �

8�I��JJJ��J��J} � �� �  �� ;i (+`�0H;8� [�� �H�H�h����� �� �� ��	  Ǐ�� �� _���  MÊ


�� ��
 �� � ��  ڐ�� ;i (+`�0� ��H�� �4  ��� � �  ��� �(+`�0� ��H��  ְ�  ְ�(+`�0H;[h�� �dZ ��ze�  �� �i �� ���hh(+`�0�;[� ��H��� �� ~�� Ȧ�� ~�� �Ȧ�� ~��hh(+`�0�;[�  ) J�� ) 


�� ) �J�� hh(+`�0�;[�  ) �� ) 




�� ) �

�� �hh(+`�0;8�	 [�� �� �d� ���  � �q�������� ⃿ ����8�� ��� �i �� ���� ��;i h(+`�0�;[� ���%�  �  �� � �	� 8� �� �i �� �ש�hh(+`�0;8�	 [�� i ���d� � ���  ���I���  � ���I��� � ���I��� � ��� � D�� e��i ��� ����� ��;i h(+`�0;8�	 [��� i$ ���� �  �  � � �  넅�i ����  � � � �  � ��� �/ �� e��i ���� �  � �  � �  �e�� � ��;i h(+`�0� ��H�� � �� � }ë(+`�0;8� [� ��H��  �� i0 �� ��  d����Y~�  ��Y~� � w�e�� ���i ���թ  ��;i h(+`�0;8� [� ��H�� �  �  ��� ��� �� �Z �z�  ��hi ����
  Ǐ� � ��� � ��
 ��  ڐ�� ;i (+`�0;8� [� �  �� �� �	��H���������� �  8��I��� x� �� �B Hh�B (�
� � 8��I��� x� �� �B Hh�B (e
�
� � 8�	�I��� x� �� �B Hh�B (e
������i �� ��L!���8�� ��� �
;i	 h(+`�0� � ⃿ �� �(+`�0� �H�H�h�  �! )���! � � )��� �$ �" �& �4 �   ���0 �(+`�0�;[� ��Y~�7���`�  �������Y~�� ��`�  ������� ��`�  �����  hh(+`�0;8� [� ��4 ک~HZ ����H� N�� ;i � � Ǐ� �� ��  �� � �� �"� ��   ڐ� ;i (+`�0� ڼ � f�z�   ְ(+`�0� �x�V ��Y �8�\ ��_ �b � �W �Z �] �` �  Ǐ�: �V � � �� �� ��   ڐx��\�J  n���\�F  n���\�B  n�� Ǐ�@ � �u\� � �~� �!� � �   ڐ(� ک~H�d\Z ���T �H� N�� ;i � � Ǐ�> � �T � � �� �-� � �   ڐ� ک~H�S\Z ���R �H� N�� ;i � � Ǐ�< � �R � � �� �'� � �   ڐ�& 0�� �  ���' 0����  ���0 0���  ���1 0��1�  ���. 0���  ���# 0��0�  ��(+`�0;8� [� �� ک~HZ ����H� N�� ;i � � Ǐ� �� ��  �� � �� �"� ��   ڐ� ;i (+`�0� x��]�J  T��y]�F  T��l]�B  T�� Ǐ�@ � �c]� � �~� �!� � �   ڐ((+`�0� � �)@��� �(+`�0�;[���]~�B �� ���]~�F �� �� ^~�J �� ��`^~�N �� �� hh(+`�0�;[���]~�B �� ���]~�F �� �� ^~�J �� ��`^~�N �� �� hh(+`�0;8� [� ��c �c �&��+�1�LB�� �R ��� �T � � �   �����] �   ��] ��L��� �F � �^~�ƥi� ���  ��   �����] �  �d�   �� ����) :��] ���[�R � �T �� � �   �����] �   �����] �  �
��   ���� ���) :��] ���i� ���  �;i (+`�0� �:  f��J  ψ�F  ψ�B  ψ�@  f��>  f��<  f��& 0�� �  ���0 0��0�  ���1 0�� �  ���. 0�� �  ���# 0�� �  ��(+`�0;8� [� �c  Ь� ���� � X� ��� � � ݱ 爢  ��i���i���  �æ pȥi���  ��� ����Ц p� �� ��� � � X�;i (+k�0�  ��(+`�0� �J  ψ�F  ψ�B  ψ�@  f�(+`�0;8�	 [�  Ь� ���� � X� ��� � �i@� ݱ�<   � ��� ����  ��  �M�� pȩ��   �� 8�
� )� � ]�� ����   ����   ��:
� )� � ]�� ���Щ���  �� pȢ   � �� ���� � X�� ;i	 (+k�0� ��H� ���(+k�0�;[� ��H�� ��i���  ��i@�  ��i��  ��� hh(+`�0� �H�H�h� ���)� ����i��  ��(+`�0� ��H�� �  ���d � �`  ���f � �i@ ��h ��  ���j �l �(+`�0� ��H��d  ְ�f  ְ�j  ְ�(+`�0� ��H��h �  �  �������  8� I��(+`�0�;[� �� �q ������ �  �� ���q �: MÊ��	 hh(+`�0H;[h�� �H�H�h� H� �d �  � �$� �i �� ���� d�� �<�~=�b�j�`~=�j�b~=<A � � U U �|��}�b�j�j�b�}�b�j�e` � � U U �~��~�a�j�b�}�a�j�`�~~ � � U U �<�~=�b�j�b�~�b�j�j�bb � � U U �|��}�b�j�b�}�b�j�j�bb � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U �<�~=�f�f�foM<�~��~~ � � U U ��<Y|9<�<�<Y<Y<�<�~=<A � � U U � � U U��~�~�~~�IU � � U U � � U U � � U U � � U U � � U U �<�~=�f�f�foM<�~��~~ � � U U ��<Y|9<�<�<Y<Y<�<�~=<A � � U U                                                                                                                                 �<�~=�b�j�`~=�j�b~=<A � � U U �|��}�b�j�j�b�}�b�j�e` � � U U �~��~�a�j�b�}�a�j�`�~~ � � U U �<�~=�b�j�b�~�b�j�j�bb � � U U �|��}�b�j�b�}�b�j�j�bb � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U � � U U �<�~=�f�f�foM<�~��~~ � � U U ��<Y|9<�<�<Y<Y<�<�~=<A � � U U � � U U��~�~�~~�IU � � U U � � U U � � U U � � U U � � U U �<�~=�f�f�foM<�~��~~ � � U U ��<Y|9<�<�<Y<Y<�<�~=<A � � U U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��""  ####    ��  ��  ��      ""``""      ��  ��  ��          ��  ��  ��                  ""``""                  ��""        ��""��""��""    ��""��""��""��""��""��""    ####            ""``""  ��      ��  ��  ��  ��  ��  ��      ��  ��  ""``      %%%%%%%%%%%%%%%eeeeeeeeeeeeeee    %"!$!&!(!*!,!.!0!2!4!6!8!:!<!>!@!B!D!F!H!J!L!N!P!R!T!V!X!e    �#!%!'!)!+!-!/!1!3!5!7!9!;!=!?!A!C!E!G!I!K!M!O!Q!S!U!W!Y!�    ������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     5               h                  Z          � �J      �    �  H z ������������������������Ѐ�������      �  d      � �                  
 �    .Fx� ` �  \��               �����           , , , , , , , ,      B �(+`�0� �H�H�h� H�Z� B[� �� �L⢥�� 	��� �  � d� ��H �̥)����� �h
 �� �� �� � �� � �� ǩ���� )�� �  D��  �� �� ��� z�h�(+@�0� ��H�� �P  ����  餭� 	�� � B �(+`�0� ��H���  ְ�� )��� � B �(+`�0) 



m� H�  ��� (+`�0H;[h�� �H�H�hH 鬅h��� )� 



m� �� �� ����� �� � �i �� ���hh(+`�0H;[h�� �H�H�hH 鬅h��� )� 



m� �� � ����� �� �� � �i �� ���hh(+`�0H;8� [�� �H�H�h� �)� � �



m� ��� �& �)� �� �� � )� ���� �i ����� hhhh(+`�0H;8� [�� �H�H�h� �)� � �



m� ���
 �& �)� �� �� � )� ����
 �i ����� hhhh(+`�0� ��H� 鬍� �(+`�0� ��H��� �(+`�0� �@� [���B �� �)����H� �)����
�d� �)�	���I�#�� �)�
���
I�#�h




͖ �#�� �� � ����� �� �� ��  X��� (+`�0;8� [� �� H�� dd�B ���� ��� �hhhh(+`�0�B � (+`�0;8� [� �� H�� dd� ���B ���@j� &j&� �����B � ��� ���;i h(+`�0�� (+`s�������0;8� [� �� H�� dd�B ���� ��� �hhhh(+`�0�B � (+`�0;8� [� �� H�� dd� ��B ���@j� &j&� �����B � ��� ���;i h(+`�0�� (+`�F�T����0� �� �@�� ����.8� �� �� �  ����������� � ���B �� � (+`�0;8�
 [� ��H�� �� ) �L
� 餩 ��  �� ��	 ���00�� �L駩  H��� :Hk�I���� E%� 9 �7� )� � �, ��� ��� �� �8�� � �	� 9 � �  X��	� E%� 9
 �7� )� � �, ��� ��� �� �8�� � �	� 9
 � �  X��	� ��  � �d� � �  � �� ����i ���L,��;i
 (+`�0� ��H��� �(+`�0�;[� ��H�� �@�   ���� �� � �i �  ������ �� �� �� �� �  �Ü� �� �� �� hh(+`�0� ��H���  ְ�(+`�0� ��H��  �;�� � �
`�~ ��� �� � �� �  La�� �   竭� ����  A��(+`�0�;[� � ڢ� ��  ��� ��� ��  �h�  ���  � hh(+` �k�0� ��H�� x�� ;� � �
 �
��  ֨��� � �� �  �� � �� �� �
`�~ ��� �� � �  �� �  �� � � � ����&�� � �
 � ��� �
 (�(+`�� � XΎ k� ;) �[i� ����� ������ � XΎ k�0�;[� ��H�� �� �>�  �� ��  谦�  �ˤ�
  :���  o��� � ְ��  � �  ת�� hh(+`� x�H��� �� � �� �  �� Κ LH��0� �� H�� �!��� �  :�� � :�� � �~�� � �� �� �(+`�0H;8� [�� ����� � �  �	����  �+��  �8�I��� :� � i�� 8�� �� B�� �� ;i (+`�0�� 8� ) ��i� �� �  � �� �  �� (+`�0H;8� [�� �
 ZHک H� {i H N�;i �� �Q��  �� �  � ��� �� �� � {i �� �  w��� �� � �  �ˊ�� �� ����� ;i (+`�0� �H�H�h� x ����	 ֨� � (�(+`�0� ��H�x�� �  W� �ڬ� �  C���l� )���� ݱ�  (�(+`�0� ��H�� x���� �
 �����
 �
�� � � � �ڬ� �  C���� )� �� ��� � � � ݱ�  (�(+`�0� ��H�� x�� �
 �����
  �(�(+`�0� ��H�� ��-� ��� �  ��  ����� ��� ���  �  � �� � ֨�(+`�0� �H�H�hx ��  � i��� (�(+`�0� ��H���� �� �(+`�0� ��H���� �� �(+`�0H;[h�� �H�H�h� )� ��� �� � )� ���i ����  �� hh(+`� ;) [(`�0� ��H��� � �(+`�0� ��H��� � �(+`�0� ��H�� �.8�  � <��~ � P�	� ���" � n� ڿ �� �� ��� �`0Od0Oh0Ol0� �� &� )� W� � � �� g�  � �Ʃ~ �  �	� �@�" ��~ � @�	� � �" ��~ � L�	� ���" ��   0��  �  ��� �(+`�0� ��H��(+`�0��;[� � �)@�t ��  ��j���  " � � �ˆ���� /ՠ0 � � �)@�( ��� ������
� �� X��� ݱ�� ݱ�I���ĥ�I� /զ �˩��  " ��hhh(+`�0� ��H� 7��  � 竀 ���  �!� 8���� �� ݱ�  �� ݱ�  � ���(+` u���d�~ �� �� (�"  �" �\	 � u���^�~ �� �� (�L��0� ��H�ڛ�  �  }�� ���(+`�0H;8� [�� �H�H�h�d 鬅�� �� 8�� ����� �����������  �^� 8��� ���� � ��� �e�� �� ������  �� � �:��� ����� �������� �






i  �� �� ;i (+`�0;8� [���Y8�  ) �P�8�  JJJJJJJ� �� )� �� �� ��.�� �ڞ� ��������ʽ� 8����� ���� ��� � ;i (+`�0� ��H�� �i JJJJJJJ Y��(+`�0H;8� [�� �H�H�h�� ����� }æ�� ;i (+`�0� ��H� ��(+`�0H;[h�� �H�H�h� �� ������� ������� �	��� ��� �hh(+`�0� ��H�� �  �������� � �i �  �����  �(+`�0� ��H��� ְ�(+`�0H;[h�� �H�H�h� )� �� ���  �� ݱ�i ����� hh(+`�0�;[� ��H�� x���  ���  � 鬦� � (�� hh(+`�0� ��H�� �  �����x���  � � � ��(�(+`�0� ��H�� �������  H� �)� ��  h��  ��(+`�0� ��H�� x �H ݱ���(�(+`�0H;[h�� �H�H�h� x�  � ���'�
 �������
  i������  ������  ���(�� �hh(+`�0H;[h�� �H�H�h� x�  � ���$�
 �������
  i�������
 ���  ���(�� �hh(+`�0� ��H��  �����(+`�0�;[� ��H� B�� ��� ��hh(+k�0� ��H��(+k�0;8� [� � �  ���� ж��� �  �0 ��� i8 �� �p  ��i� �� �  � ���  �  �¦� � hhhh(+`�0�;[� ��  � ���  竦 ӳ�� ���hh(+`�0� � ���� ��  � �%� ��  � � � ���  � � �� �� (+`�0� ڼ  � ��� ְ(+`�0H;8� [�� �H�H�hH)��h)������ �  ����� �  ����� �  ����������� ���� � � ��8��
 �JJ� �  =��� �i �� ��ή���� �  ���  ��� �i �� �� �i �� �� �i �� �� �i �� � 8�

�	 
�
 �� � �i ��Щ�� hhhh(+`�0� ��H��� ְ�� ְ�� ְ�(+`�0��;[� ��
 �� )� 

m��� )� �� i �� �� i ��
� �� L�� � )


H� )
�� )��  )�� � � � � � �  ���I�  )�� )��)���h��

��H�I���JJ� ) m��� � %� hhhh(+`�0H;[h�� ���J�� �i �� �� 8� �� �� � �� ��%���� �i �� �� 8� �� �� � ����  h(+`�0H;[h�� ���J�� �i �� �  8� �� �� � �� ��%���� �i �� �  8� �� �� � ����  h(+`�0H;[h�� �H�H�h����� ��  �8�� �� �,� q��  �"�� �� ���  �� �� �������hh(+`�0� ��H�� ���� � �
 )� 

m��� �� �(+`�0���� � � �
 )� 

m��� �� (+`�0�;[� ��H���� _��� ���Z�   _�z�����h(+`�0� ��H� =��(+`�0H;[h�� �H�H�h� �� ���JJ�  � ���������h(+`�0� ��H����(��� Ǐ�  ��� � ��� � � �
 �  ڐ�(+`�0;8� [� �  ���  �n����� �  �î��  �ڼ  �
 ) H



e��	 H



m��� ��  �  �������hm��he�� � � � ��i ��Э� ְ;i (+`�0;8� [� ��H����W��� �  ���  �G�� �  ����
 JJe���  i ����� ��ʩ����  ���8��	 ��� ְ @��� ;i (+`�0�;[� ��H��  z��� ��� hh(+k�0� ��H��(+k�0;8�
 [�  �� �  ���� ��ک~���Q ��� ���� ��	�dd�	 ж�� � ���(`~�i�� �(`~� )� �i` � ��	��  ��� ��Ħ� ;i
 (+`�0�;[� �� !��� � 竀�hh(+`�0;8� [�� � ��  �ª�� i �� �  � ��	 ��:`~)� ��  � �H� ��h������� hhhh(+`�0;8� [�I �  ����  Ǐ��
 �  � � � � �~� �  ڐ�  Ǐ�i �
 � 0� � � � �~�  ڐ�  ��ک~��PQ ��� ��

	 � � ��  mǆ� �� ��  I �  I ������i  ���ݠ@�!�  ����� pȩ  0�����  ���  0��  �  ��;i (+`�0� ��H�� � �   ����� � ��  �i  ����(+`�0� ��H��� ְ�(+`�0� �H�H�h� ) 




m��� � �<  ��i  ����  ��  �(+`�0� ��H�� � ��  �(+`�0�;[� ��H�� ��  Ǐ�  � �� �8��J� H�
 ��  ڐhJJJJ��hh(+`�0�;[� ��H�� ��  Ǐ�  � �� �8��J� H�
 �� ���  �;�  ڐ��  � hJJJJ��hh(+`�0H;8� [�� �H�H�h����� )� JJJe��) ��  ��  �������;i (+`  �                            �0�;[� ��H�� ��  Ǐ�  � �鼝 �8��J� H�
 �~�  ڐhJJJJ��hh(+`�0H;8� [�� �H�H�h� ��)� ���)� 8��!���e��  �� �  �������  �;i (+`�0H;8� [�� �H�H�h� ��)� ���)� �8��!���e��  ��ʽ  � �����  �;i (+     ,�    PR�s     ,|          �joV�EH9�$  �{w�^sR�f�V.F�9)�0�A��$E�$�b"�f�V.F�9)�0�R|F�5�H�w_vJ�AL9�$�$E�0  �`?w�^0J�=I-�   �E�,D� �jqR�A�1%  ��|��g�o�G�c���@sf1^�Im-+%��9a$b�"�-@M M N�M�@�|��o
`-�9chs@5`5�9BCJ�V�c�t�3��>�)��C��>�)��CUU�yQ�)�>�T�R$9Gb�{%��UU�t��U.W�6�W�8]]_vS`9�{UU�� z5]>�::WCr�-�6�[8U�z�UU�<>BO�k�!�>�W�i�rw9��'<�  !�-�6�C�{:�K�1L>v_-A�U�f�G�{��F�>w>42�%�*�����~G}�\k-��,MA6f>�!�6�K�1�>�;�C	�_�                                ����H����(+`                                �����>`~)� ��	���m���  � �(�(+`�0� ��H�� ��x���  ��(�(+`�0� ��H�� ��x8��� ��� � � ��(�(+`�0� ��H�� �  ��� )� �m������ )� �m������(+`�0;8� [� ��H�� � !��  ���� )� �(m��H�  )� �� � ���>`~�����z� �Р�� )� �(m��H�  )� �� � ���>`~�����z� �Ы� hhhh(+`�0�;[� ��H�� ������ )� �<m��H�  )� �� � ���>`~�������� H�>`~)� �h�� z� ����� )� �Jm��H���	���  ���  )� �� � ���>`~�������� H�>`~)� �h�� z� �����	���  ���������� hh(+`�0� ��H�� ���� ��� �����8�����(+`�0H;8� [�� �H�H�h� )� �� �:�� e�8� I�����J���� [�%����� �hhhh(+`�0;8� [� ��H�� ���$u���� ��� �)@�I@�
�	 �J���J�� ��J� �  ����� �����   ������г���hhhh(+`�0) �� �  �
����(+`�0�� 
������ ��:(+`�0� �  �4�  �� �� ���:� �" �ÀH�)�h��H��h� �  �興��� (+`�0H;8� [��  �LE�� �D�:�� �T������k���~H� ��H� � H� {i  H� � �xk(���٫� �'� �H� �  �  � ��h:�J��  �  �������;i (+`�0;8� [� �� H�� ��l� �H:�� �T������k��
���~H� ���H� � H� {i  H� � �xk�(����� ��  � �� ��
� �:�J���
������� hhhh(+`�0H;8� [��  �Lz�� �N�:�� �D������`�� �e�� � �e�� �� �6�H{i  H� � �x`�(����� �5��e��e��� �ʈ� �  �  � �:�J��ʈ��  �  ���;i (+`�0H;8� [��
�/e�ej)�����  �������e�����e�٠  � hhhh(+`�0H;8� [�� �H�H�h� ����  � �Ŋ8�J8��c�c�FU��_��>�)��C��>�)��CUU���<1!�-�B�df�Ip^0s�|�UU�t��U.W�6�W�8]]_vS`9�{UU�� z5]>�::WCr�-�6�[8U�z�UU��>�)��C��R�1�QR��R�1�QR  ,��S��f{�z�Uv�~/~�	��5�� ��5�R�yZr�~]5�.^7�_��� ��5�R�yZr�~]5�.^7�_�    �� �� �� �� ��� ��� ��� ��� �� �� �� �� ��� ��� ��� ��� �� �� �� �� ��� ��� ��� ���  �� � � ��  0H;8� [�� �H�H�h� � ǅ� �)� � �� �����  ک  ��� ��� � � h�� � JJJ�)�� �զ�  

��)��JJ)�i 0���  ���
i 0��      �
"�� � @      �
��  @      �
��  @�     �
 ��@��6       
 3!@ �       
 25@ ��      
 @ �  
    
 -6@��  
    
 	4@��  
    
 "@�  
    
 '@��      
 #?@��      
 2H@�       
  c@�      
  G@ ��  
    
 7L@ ��      
 3X@ ��  
    
 5@��  
    
 Z@�       
 
X@��      
 *d@�       
 d@�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �:	��  ���  竀�(+`�0� ��H�� ��  ����(+`�0� ��H�� ְ�(+`�0H;[h�� �H�H�h��  �x�  �� �i �� ���  �
�� ��  (�h(+`�0� ��H��  �(+`�0H;[h�� �H�H�h��  �x�� ������       ������������������������������������V�����������������������`������������ �@����              *              H���  �(+`�0�;[� ���� �� ��� �  X����  hh(+`�0�;[� ��H��� ��7! �=! �=! ��ް�  �� �� � ���i �� ��ѥ�^D ^D �  [� ��H�� ��.�8�  I��

m��  )� � �� � ���i ����� hh(+`�0� ��H�� � +��  � ��  ߇                                                                                                                                                 ^D ^D �  [� ��H�� ��.�8�  I��

m��  )� � �� � ���i ����� hh(+`�0� ��H�� � +��  � ��  ߇                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �   f�  �   Z���  0�� ��� H ��h���(+`�0� �_�~ ����� �� �� �L�ҭ��  �� �����  �-� �� �� " â� �� �` ݱ ��� X�� �� �J ��� �C�   �͢  �� �3��  �,� �� �� " � �� �����^�~ ���(+`�0�O��" "�_�#^NIB2�-�-�-e!��O����_�#^NIB2�-�-�-e!��O����_�#^OIB2�-�-�-e!��O����_�#^PJB2�-�-�-e!��O����_�#^PJB2�-�-�-e!��O����_�#^QKB2�-�-�-e!��O�`��_�#^RKB2�-�-�-e!��O�`��_�#^RLB2�-�-�-e!��Oi`��_�#^SLB2�-�-�-e!��Oi@��_y#^TMB2�-�-�-e!��OI@��_x#^TMB2�-�-�-e!��OI@��_x#^UNB2�-�-�-e!��OI ��_W#^VNB2�-�-�-e!��O) ��_W#^VOB2�-�-�-e!��O) ��_V#^WOB2�-�-�-e!��O) ��_V#^XPB2�-�-�-e!��, �� ���� �� И��	� ��� �ѭ��  р� ����	 ��� �� ��hh(+`�0� �H�H�h� ��� pȫ(+`�0� ��H�� �� �  "  � ЬH ��h X��
��  竀�
��  Ǐ�
i � � � � ��
 �� �  ڐ�  竀˫(+k�0� ��H��(+k�0� ��H�� �   ���,�(+`�0� ��H��, ְ�(+`�0H;8� [�� �H�H�h��JJJJ�d� ���,J�F���  �������  ���� �e�� ��ܩ�������  ����� �8�,� �� �;i h(+`�0H;[h�� �H�H�h� )� m,�� � ��  �,�  ��  ����h(+`�0� ��H�� �) ��JJm,��  �(+`UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUF  |�s    |�s                  ���%�B� �_~e�<*�%O���6x**�%O��O��3'�&�&*�f��\G�:X.�-n!��.&�R��&*� ��\G�:X.�-n!��.&�R�2*�)N! ��Z[�J�F:�-)�f�i\=R'�&�&*�F�����[ko�4_~e�<��&�&*�f����[���.����&���@���I V`b�j��c�c�FU��_��>�)��C��>�)��CUU�yQ�)�>�T�R$9Gb�{%��UU�t��U.W�6�W�8]]_vS`9�{UU�� z5]>�::WCr�-�6�[8U�z�UUm �_�mz�~N��L!6�F[g�  ,��S��f{�z�Uv�~/~�	��5�� ��5�R�yZr�~]5�.^7�_��� ��5�R�yZr�~]5�.^7�_� U�              #\\     � � � �2 @&     �      �               //  �               
     3  �5`     ��7@0�X@ @@  � D2 �#   ���3� �#� �# �#                                �       ��  ��D1�F1� H1��J1��L1��N1��`1@�b���d�    "  6�  �WYX               ��   �                 �              �X                                                      i  � E   I         O           )   �� P         �                        O              ��   M        P   �      X :   $                            @     �  �                        �                        @0   0�   ��7@0�X@ @@ ��  h  �%                                                                                                           B                                                                          xc         �Xxcxcxcxcxcxcxcxcxcxcxcxcxcxcxc                �                                           ��                                                         �    �                     X :   $                             @     �  �                        �                        @0   0 @  ��7@0�X@ @@  �  �  �'                                                                                                           b                                                                          xc         �Xxcxcxcxcxcxcxcxcxcxcxcxcxcxcxc                �                                           ��                                                         �    �                    �T              ��         �  r @       �0       @��6    �          wY                   �:   0``\6
��:�:�T@ @  ��  �r @*    �@z��B:                                                                                                � �                                                                         �T                                                          �                                           ��                                                         �                        e�        �   ��      � � �  D E    � �@     @�            D   W�               	  <T�20�G����4J<T�EE5 �  �D h,   �h<��j<l<�n<��,
�l���,
��l �l�l         �       ��  � �(� �(�  )��9�9� 9 9�
99�9� �                            ����  �                                �

J � �  � �>                                            < <       �   c          �       � 5         �                                       K � KL     �             ��           !��      @ p �   E     �      @�            /  �Q	            ,�    <T�20�G  ��4J<T�EE5 �   	 �.   ���~���~��~��~��>
�~���>
��~ �~�~         �       � �  �  9� "9� $9��&9�(9� *9 ,9�.9@9�B9� �                            ��
   �                                �
J 0@ p  � �>                                           & <       �   c          �       � 5  �      �                                       K2� KL                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �n �nZ�� �Z�����Z���Z�� :� z��f��bZ��bZ��`Z�.Z��,Z��LZ��NZ                                                                                                                                                                                                                                                                                                                          >  $>@ (>` ,>�  ~� $~� (~ � � �$�@�(�`�,��� ���$���(�                                                                       ��L���L��L                                                                                                                   ��                                                                                                                            �� _ � ��_ ������ ���_                                                                                               �� _ � ��_ �                                                                                                               �� _ � ��_ �                                                                                                               ���������������������������������������������������������������Ɠ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� W �������������                                                                                                                                                                                                                                                                                                                                                      W �������������                                                                                                                                     �������������������������Z�Y�44�����(#O%!"3����5) �������������������������Z�Y<�)"jkkl>>M%L>>>>	�������������������������Z�Y�S�4������E9)*+3����������������������������������������������������������������<Z�Y;�;�����������������������������������������������������������������������������������Z�Y�������U?	
+C�����5)�������������������������Z�Y<�^)joooZ=%!">1$L>>>	�������������������������Z�Y�S���������4::�����������������������������������������������������������������NZ�Y;�;�����������������������������������������������������������������������������������Z�Y�������5 $/+3������E��Z�Y<�$N%LYoooZM/L>>"O/L>>	**��Z�Y�S�������TU	S�����������������������������������������<Z�Y;�;������������������������������������������������������������Z�Y��������5 !"+3�������E	+��;Z�Y<�$"	YoooZ %">>>LO/L>>+ ��Z�Y�C�����E	
S��������������������������������������<<<<<<<<<<<<<<<<<<<<<<<<��;<Z�Y;�;������������������������������������������������������������Z�Y���������5	
+3�������TU #��;Z�Y<�%?N	1zoooZ/L>>>LO/L>	 "��Z�Y�S�����US�������������������������������������<<<<<<<<���������    ����<Z�Y;�;�����������������������������������������������������������     ��Z�Y���������E)+3�������U	
+����  ��;Z�Y</�/??",YooZ/L>>" #O%"	
<<<<<<<<<<<<<<<<<� �  ��Z�Y��C����5)**S������������������������������������ ��<Z�Y;��;����������������������������������������������������������;;;;;;;;;<;<;<;<�$/�Z�Y����������53�������U	 "#"#$����;;<;<]^�Y<��1"	?zoo|,>>L%"	$2323���/]cd�Y��S�����4:5C�����������������������������������""""""""##"#"#"#$�@DB��l;</]cd��Y;m���;<����������������������������������������������������������2222222233232323���@DDD���/]cd���Y������������������E	M��FDDDB�.;<;<]cd����Y;</�.;1	,z|,">>,O/L	�FDDH���/cd�����Y���S�����4US�����������������������������������;<;<;<�� .;<;<;<cd������Y;<m����;<;<;<;<;<;<;<;�����������������������������������������������������������/��� .]cd�URRRS�Y�����������.�������������������U<;<;<;<;<;<;<��� ]bbbbbbcd�UV��Z�Y;<�����lml%"?",�>>MO/L��]cfffffffffg�UV��Z�Y����C�US�E	C�����������������������������������������ǔ������/]cd����������UV�Z�Y;<m����l���������������������������������������������������������������/]cd�URRRRRRRRRV�Z�Y�������������������U	+�������./]cd�UV      <Z�Y;<��.lml%"	1",�,!u"O/L���������]cd�UV��Z�Y��S�53�UC���������������������������������������� ]cd�UV�Z�[;<;m�;������������������������������������������������������������� �]cd�UV WX`a]������UST���������U	** #��� �]cd�UV <WX`a];</�l/"	,>>,-u��>OL�� ]cd�UV����������������WX`a/��ST�E	S����������������������������������;</��]cd�UV <;<;<;<;<;<;<;</WX`a\����;������������������������������������������������������������]cd�UV./WX`a\��.��U	
ST������E	+35)*#m]cd�UV ;<"#"#$WX`a\��.;<;<;<;<;<;<;<;<"	?L>>>>,u>> )ld�UV�!$23234WX`abb  bbbbbbbbbbbbb
SUST��������������������������������<<<<<<<<<<Z��Y1!"#"#"#"#$WXeff  fffffffffffffff����������������������������������������������������������Z��Y123232323WX��  ����������������U	
S�����E+3��45)#m/Z��Y<<<<<<;<;<����;<;<;<;\WRR  RRRRRRRRRRRRRRR	>">>M%L�Z��Y�������;<;<�  ���


S�������������������������������<<<<<<<<<<�Z��Y;<;<;<����������;<;<;<@DDB���������������������������������������������������������������Z��Y�/�����������lmlmlm/�/DDDH��l�5S����E)+3�����5) _m�Z��Y�;</�����������.���.;<;<�DDE����%"+"� ">>>>/L�Z��Y���������������;<;<;<ʻ���/��FGH���lC������������������������������<<<<<<<<<<�    ���./����lm��������������������������������������������������������������������������������    ���������--������lm�����lmlm�l�E)C����5)+3�������5),}~~�����=>?O�������%1"	"�>>>�>>>>MLZ��Ylmlmlm�IJKL���lml;<;<;<��llmlmlml+C������������������������������<<<<<<<<<<Z��Y��������/����������������������������������������������������������Z��Y;<<<<<mlmlmlmlml;;;;;<���l��5)3������53���������5)**Z��Y/�lm%%$	11L>>>>>>>>>>,)Z��Y;;;;;;;;;;;;;;;;;;;;<�;<;3�������������������������������<<<<<<<<<<Z��Y/�l���������������������������������������������������������������������Z��Y;<<<<<<<<<<<<<<<<<<<� ������MN��MN����������� �!�>v n�}C_� l�>��|�!�w u:�?� FO?^h�>nnZ��Y��l<   ��������������������r�?�(2.z?� ��z�>�+��p , UzH� �9�� 8 ��?4 UZ��Y<<<<<<<<<<<<<<<<;</�������������������2 [ xn?���'�9� � ��>+6l�T ��=] ��>�?� (Z��Y�l;<;<;<"#��������7vl>��@1 � 0 �'�� ?   @   v>5 g=_�$�� �**� V <<<<<<<<<<<<<<<<<<<<<<<<<<<;<;<		!"#$23!!"#O _
a?- 'l}D�. ��=g ��~�?Zc� �3 � �U�>{��^$�� 

�;<;<;<23!$123!i n & 0~��u �7 ; IC�E   	   d3?� 	D<  m�
.
��!"##"$4;<MN�1!"#"#"#"n h]��� ��?� I/>� {0l@A� �a�?c&� ] �,1� /
��.	
���2332  MN12323232)
� - HOQ�s �$�#� � �4�AT �%�$� � t5>R }�[f'<� Z�Y;</���	���
lmlmlmlm����;</�� )  h%�� 3 �
�?K 4�F�a �W�^e ��=� K��� � Z�Y
bbb\��	�/��!� � !�  �:U?� �?� ��>� q	 o 
�S b H
� S Z�Y;<lfffm��lmlmlmlm/����1!"#"#"#"#"�W'�;u7�4m �}	G V �D$	�Z �72'� N�!M�4 T Z�YZ���Y������232323232l � F �� � ��R0 Z{0rO�L�  ,�4> �tf � Z�Y;Z��UVlml<;<;<;</�����.�&4F� ��
�`� 6 0!��w%y��S f R&m�� <Z�YZ��Y������ .;��A���+ ��3' y.Xk < 8l � �	v� ?�i� a Z�Y<WRRV�l����.;<:�f'vD�6�
/(�x
n&�n�  �@ �  GZ�Y���#"#"#"#"��MN;<;<;b RJRJ    J v     �t     �     � (     �      4 �Z�Y;<;<;<�;<;<;<32323232!#"��������53:US�����������������������5<Z�Y132��!"#"#"#"#"#"#"?%L>	
	M%	/]^�Y���232323232323S������������������������������<]cdUV"#"#"#"#"#"#"#@DB  ����������������������������������������������������������/ldUV23232323232323;<;<DDDDB ;�������U34:�����������������������E)**<;<Z�Y@DDDDDDD 1$)+"	
,%"Z�Y<;<�;<;<;<DDDDDDDH S�����������������������������</��Z�Y�@DDDH/.�������v�����������������������������������������������������   �.;<;<;<;<;<DDDH/�� ;�������4�E3������������������������5) m/���   ��./.@DDD/]bbb\� 1$)*+=	��	����}~�������./��;<;<;<;<;<;<;<DDDH�lfffmlC����������������������������<����Z�Y�������������/������.FGH�^���Y�������������������������������������������������������������Z�Y������������lmlmlmlmlm���/ld���Yl������������������������������������5)+#m���Z�Y��������Z����Y.11$N)*="

	���Z�Ylmlm������llmlmlmlmlmWRRRRVl+3�����������������������������m	�Z�Y�������������������������������������������������������������	��Z�Y;mlmlmlmlml<;<;<;<<<<<<<<<mlmlml�������������������������������������5)**M_m	�Z�Y$)=>��Z�Y�;<;<;<;<;<;<;<;<;<;<@DDB;<;;;;;;;;;;;;**+3������������������������������<;<��Z�Y����.FDDDB����������������������������������������������������������/��   ���������.�������FDHl��������������������������������������445*****,m����   �lmlmlm����lmlmlm��������^N###%L)*)}~�����������;;;;;;;;;;;;+344�������������������������������mlZ�[\�;mlmlmlmlm���������������������������������������������������������������WX`a\.���l����������������������������������������E)*+34445)*,WX`a\;<;<m�$%^�)1L)**WX`a\./��;+3����������������������������������WX`a\.;<;<������������������������������������������������������������WX`a\.���l�����������������������������������������534�����45)WX`a\;<;<��$2N#O$N),)WX`a\.��l*+C����������������������������������WX`a\.;<;<������������������������������������������������������������WX`a\.��;���������������������������������������������������5)WX`a\;<;<��^#2#O_%?L,!!^)WX`a\.��*+)34�����������������������������������WX`a\.;<����������������������������������������������������������������������������������������445�,"3���������������������������������������������������������������������������������5)***M_%!"35,%$$LC���5%?$N######%1$###2##%1L�	�,)ff,-.,N#---.	
I>fjl#	+345+C����������������������������������������������������v�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E)***
=f=<g<<gf=>	*+3US�����������������������������������������������������������������������������������5)*�34����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������45)+35)*


=fg=>	
+34U	C�����������������������������������������������������������������������������������5)+)*C������������������������������������������������������������������������������������������������������[[[[[[[[[[[[[[[[[[[[[[[[    \[\[\[\[\[\[Z��� Y\[\h   Y\[\[\[\[\[\[\[\[����������������������������������������������������������[[[[[[[[[[[[[[[[[[[[[[[[    lklklklklklkj��� ilkl    ilklklklklklklklk




CU[[[[[[[[[[[[[[[[[[[[[[[[    [\[\[\[\[\[\h��� g[\[Z   g[\[\[\[\[\[\[\[\����������������������������������������������������������[[[[[[[[[[[[[[[[[[[[[[[[    klklklklklkl ���  klkj    klklklklklklklkl����������������������������������������������������������[[[[[[[[[[[[[[[[[[[[[[[[    \[\[\[\[\[\[Z��� Y\[\h   Yg[\[\[\[\[\[\[\[����������������������������������������������������������[[[[[[[[[[[[[[[[[[[[[[[[    lklklklklklkj��� ilkl    ilklklklklklklklk9[[[[[[[[[[[[[[[[[[[[[[[[    [\[\[\[\[\[\h��� g[\[Z   g[g[g[\[\[\[g[\[\����������������������������������������������������������[[[[[[[[[[[[[[[[[[[[[[[[    klklklklklkl ���  klkj    klklklklklklklkl����������������������������������������������������������[[[[[[[[[[[[[[[[[[[[[[[[    \[\[\[\[\[\[Z��� Y\[\h   Yg[\[\[\[\[\[\[\[����������������������������������������������������������[[[[[[[[[[[[[[[[[[[[[[[[    lklklklklklkj��� ilkl    ilklklklklklklklk9	[[[[[[[[[[[[[[[[[[[[[[[[    Y\[\[\[\[\[\h��� g[\[Z   g[g[g[\[\[\[g[\[\����������������������������������������������������������[[[[[[[[[[[[[[[[[[[[[[[[    ilklklklklkl ���  klkj    klklklklklklklkl����������������������������������������������������������[[[[[[[[[\[\[\[\[\[\[\[Z    g[\[\[\[\[\[Z��� Y\[\h   Yg[\[\[\[\[\[\[\[����������������������������������������������������������[[[[[[[[klklklklklklklkj     klklklklklkj��� ilkl    ilklklklklklklklk+9)[[[[[[[[\[\[\[\[\[\[\[gh    Y\[\[\[\[\[\h��� g[\[Z   g[g[g[\[\[\[g[\[\����������������������������������������������������������[[[[[[[[lklklklklklklkl     ilklklklklkl ���  klkj    klklklklklklklkl����������������������������������������������������������[[[[[[[[[\[\[\[\[\[\[\[Z    g[\[\[\[\[\[Z��� Y\[\h   Y\[\[\[\[\[\[\[\[����������������������������������������������������������[[[[[[[[klklklklklklklkj     klklklklklkj��� ilkl    ilklklklklklklklkS5[[[[[[[[    Y\[\[\[\[\[\h��� g[\[Z   g[\[\[\[\[\[\[\[\����������������������������������������������������������[[[[[[[[ZYZYZYZYZ       ilklklklklkl ���  klkj    klklklklklklklkl����������������������������������������������������������[[[[[[[[jijijijij      g[\[\[\[\[\[Z��� Y\[\h   Y\[\[\[\[\[\[\[\[����������������������������������������������������������[[[[[[[[[\[\[\[\h          klklklklklkj��� ilkl    ilklklklklklklklk
S[[[[[[[[klklklkl         Y\[\[\[\[\[\h��� g[\[Z   g[\[\[\[\[\[\[\[\����������������������������������������������������������[[[[[[[[ghghghgh           ilklklklklkl ���  klkj    klklklklklklklkl����������������������������������������������������������[[[[[[[[                    g[\[\[\[\h\h ��� Y\[\h   Y\[\[\[\[\[\[\[\[����������������������������������������������������������klklklkl                     klklklkl    ��� ilkl    ilklklklklklklklk\[\[\[\[Z                   Y\[\[\[\h   ���� g[\[Z   g[\[\[\[\[\[\[\[\����������������������������������������������������������lklklklkj             T�U   ilklklkl   �����  klkj    klklklklklklklkl����������������������������������������������������������[\[\[\[\[ZYZYZYZ     T���   g[\[\[\h  ������ Y\[\h    g[\[\[\[\[\[\[\[����������������������������������������������������������klklklklkjijijij     W����   klklkl  ������� ilkl      klklklklklklklk\[\[\[\[\[\[\hgh      W���   ghghgh �������� g[\[Z   ]^ghghghghghghghg����������������������������������������������������������lklklklklklkl              e       ���������  klkj   mn               ����������������������������������������������������������hghghghghghgh]^           d     ���������� Y\[\h       YZYZYZYZYZYZY����������������������������������������������������������             mn     d          �����   ��� ilkl        ijijijijijiji                       �������������� YZ ��� g[\[Z      Y\[\[\[\[\[\[\����������������������������������������������������������                      ��������������  ij ���  klkj      ilklklklklklkl����������������������������������������������������������YZYZYZYZ             ��������������YZY\h��� Y\[\h   YZY\[\[\[\[\[\[g[����������������������������������������������������������ijijijij            �����    ijil  ��� ilkl    ijilklklklklklklk\[\[\[\[Z          �����YZYZYZYZYZY\[\[Z ��� ghg[Z   g[g[g[\[\[\[\[g[\����������������������������������������������������������lklklklkj       d ����� ijijijijijilklkj ���    kj    klklklklklklklkl����������������������������������������������������������[\[\[\[\[Z    e  �����Y\[\[\[\[\[\[\[\h ����   gh   Y\[\[\[\[g[g[\[\[����������������������������������������������������������klklklklkj   e  ����� ilklklklklklklkl   ����       ilklklklklklklklk*+\[\[\[\[\h   d �����YZY\hghghghghghghgh    ����      g[\[g[\[\[\[\[g[\����������������������������������������������������������lklklklkl     �����ijil                    ����      klklklklklklklkl����������������������������������������������������������[\[\[\[\[Z   ����� Y\[\h             YZYZYZYZ����     ghghghghghghghgh����������������������������������������������������������klklklklkj  ����� ilkl              ijijijij ����                    +3:\[\[\[\[\h �����YZY\[\[ZYZ          Y\[\[\[\[Z ����  pq               ����������������������������������������������������������lklklklkl  ���� ijilklkjij    YZYZ  ilklklklkj  ��������������������������������������������������������������������������������[\[\[\[\[Z ����Y\[\[\hghgh    ijij  ghghghg[\[ZYZ�������������������������������������������������������������������������������klklklklkj ����ilklklRS    ghgh         klkjij ��������������������9	\[\[\[\[\h ����ghg[\hbc                   g[\[\h  de                 ����������������������������������������������������������lklklklkl  ����   kj  01223       YZYZYZ    klkl T���    YZYZYZYZYZYZY����������������������������������������������������������[\[\[\[\[Z ����]^egh  @AB>CD      ijijij    ghgh ����    ijijijijijiji����������������������������������������������������������klklklklkj ����mn     :=B7L;      g[\[\h]^       ���    Y\[\[\[\[\[\[\9)\[\[\[\[\h ����      @<ANBABD      klkl mn    ���    ilklklklklklkl����������������������������������������������������������lklklklkl  tuuv      5LBABLN9     Y\[\[Z     YZYZ      Y\[\[\[\[\[\[\[����������������������������������������������������������[\[\[\[\[Z ����      JFGHHGHK     ilklkj     ijij      ilklklklklklklk����������������������������������������������������������klklklklkj ����YZYZYZ          YZY\[\hgh  YZY\[\[ZYZYZY\[\[\[\[\[\[\[\+9	\[\[\[\[\h ����ijijij          ijilkl     ijilklkjijijilklklklklklklkl����������������������������������������������������������lklklklkl  ����g[\[\[ZYZYZYZYZY\[\[\h  Y\[\[\[\[\[\[\[\[\[\[\[\[\[\[����������������������������������������������������������[\[\[\[\[Z ���� klklkjijijijijilklkl   YZilklklklklklklklklklklklklklk����������������������������������������������������������klklklklkj ����Y\hghg[\[\[\[\[\[\[\h   ijghg[\[\[\[\[\[\[\[\[\[\[\[\[\3U\[\[\[\[\h ����ilklklklklklklklklkl   Y\[Z  klklklklklklklklklklklklkl����������������������������������������������������������lklklklkl  ����g[\[\[\[\[\[\[\[\[\h   ilkjghgh����������������������������������������������������������[\[\[\[\[Z ���� klklklklklklklklkl   Y\[\h d  YZYZ                                                                              klklklklkj ����Y\[\[\[\[\[\[\[\hgh   ilkl  deeijij                                                                              \[\[\[\[\[Z����ilklklklklklklkl     Y\[\[Z    ghgh                                                                              lklklklklklklklklklk[\[\[\hghgh     ilklkj            YZ  YZ                                                                    [\[\[\[\[\[\[\[\[\[\klklkl          ghghgh            ij  ijYZ                                                                  klklklklklklklklklkl\[\[\[Z                         YZgh  ghij                                                                  \[\[\[\[\[\[\[\[\[\[lklklkj                         ij      gh  YZYZYZ                                                          lklklklklklklklklklkl\[\[\h         YZYZYZYZ        gh    dd    ijijij                                                          [\[\[\[\[\[\[\[\[\[\[lklkl          ijijijij                   Y\[\[\[                                                          klklklklklkjij  ���Y\[\[\h         Y\[\[\[\[ZYZYZYZ            ilklklk                                                          \[\[\[\[\[\[\[Z ���ilklkl �����    ilklklklkjijijij           Y\[\[\[\                                                          lklklklklklklkj ���g[\[\[Z����� YZY\[\[\[\[\hghghgh         YZilklklkl                                                          [\[\[\[\[\[\[\h ��� klklkj����� ijilklklklkl                ijg[\[\[\[                                                          klklklklklklkl  ���Y\[\[\h���� Y\[\[\[\[\[\[Z            e  gh klklklk                                                          \[\[\[\[\[\[\[Z ���ilklkl ���� ilklklklklklkj                  ghghghg                                                          lklklklklklklkj ���g[\hgh      ghghg[\[\[\[\[ZYZYZYZ   wx                                                                       [\[\[\[\[\[\[\h ��� kl              klklklklkjijijij   yz                                                                       klklklklklklkl  ���Y\[Z            Y\[\[\[\[\[\[\[\[Z  yz    YZYZYZYZY                                                          \[\[\[\[\[\[\h  ���ilkl            ilklklklklklklklkj  ��    ijijijiji                                                          lklklklklklkl  ����g[\[ZYZYZ  YZYZY\[\[\[\[\[\[\[\hghT�U  ee g[\[\[\[\                                                          [\[\[\[\[\hgh ����  klkjijij  ijijilklklklklklklkl   ����U  e klklklkl                                                          klklklklkl    ���  Y\[\[\hgh  g[\[\[\[\[\[\[\[\hghT������� d Y\[\[\[\[                                                          \[\[\[\[\h    ���  ilklkl  RS  klklklklklklklkl   �������X  dilklklklk                                                          lklklklkl     ��� ghghghRSbc  g[\[\[\[\[\[\[\h  T���X       g[\[\[\[\                                                          [\[\[\[\[Z    tuv        bc   RSklklklklklklkl   ���X       d klklklkl                                                          klklklklkj    ���             bcghghghghghghgh  T���        dY\[\[\[\[                                                          \[\[\[\[\h    ���                               ���X  �����  ilklklklk                                                          lklklklkl     ���              YZYZYZYZYZ      W�X   ����� Y\[\[\[\[\                                                          [\[\[\[\[Z    ���              ijijijijij           ������ ilklklklkl                                                          klklklklkj    ���YZYZ          Y\[\[\[\[\[ZYZYZYZYZYZ������Y\[\[\[\[\[                                                          \[\[\[\[\[Z   ���ijij        ilklklklklkjijijijijij������ilklklklklk                                                          lklklklklkj   ���g[\[ZYZYZYZYZY\[\[\[\hghghg[\[\[\[\[ZYZYZY\[\[\[\[\[\                                                          [\[\[\[\[\[Z  ��� klkjijijijijilklklkl      klklklklkjijijilklklklklkl                                                          klklklklklkj  ��� ghghghghghghghghghgh      ghg[\[\[\[\[\[\[\[\[\[\[\[                                                          \[\[\[\[\hgh  ���                     T��U    klklklklklklklklklklklk                                                          lklklklkl     ���                    W���U  Y\[\[\[\[\[\[\[\[\[\[\[\                                                          [\[\[\[\[Z    tuv  YZYZYZ      YZYZYZ    ��X]^ilklklklklklklklklklklkl                                                          klklklklkj    ���  ijijij      ijijij       mng[\[\[\[\[\[\[\[\[\[\[\[                                                          \[\[\[\[\[ZYZ ���g[\[\[ZYZYZY\[\[\[ZYZ       klklklklklklklklklklklk                                                          lklklklklkjij ���  klklkjijijilklklkjij      Y\[\[\[\[\[\[\[\[\[\[\[\                                                          [\[\[\[\[\[\[Z����  ghg[\[\[\[\[\[\[\[\[Z     ilklklklklklklklklklklkl                                                          klklklklklklkj ����    klklklklklklklklkj     g[\[\[\[\[\[\[\[\[\[\[\[                                                          \[\[\[\[\[\[\[Z ����   g[\[\[\[\[\[\[\[\h      klklklklklklklklklklklk                                                          lklklklklklklkj  ����   klklklklklklklkl      Y\[\[\[\[\[\[\[\[\[\[\[\                                                          [\[\[\[\[\[\[\[ZYZ����  ghg[\[\[\[\[\[\[Z     ilklklklklklklklklklklkl                                                          klklklklklklklkjij ����    klklklklklklkj    Y\[\[\[\[\[\[\[\[\[\[\[\[                                                          \[\[\[\[\[\[\[\[\[Z ����   g[\[\[\[\[\[\h    ilklklklklklklklklklklklk                                                          lklklklklklklklklkj  ����   klklklklklkl     g[\[\[\[\[\[\[\[\[\[\[\[\                                                          [\[\[\[\[\[\[\[\[\[ZYZ����  ghg[\[\[\[\[Z     ilklklklklklklklklklklkl                                                          klklklklklklklklklkjij ����    klklklklkj    Y\[\[\[\[\[\[\[\[\[\[\[\[                                                          \[\[\[\[\[\[\[\[\[\[\[Z ����   g[\[\[\[\h    ilklklklklklklklklklklklk                                                          lklklklklklklklklklklkj  ����   klklklkl     g[\[\[\[\[\[\[\[\[\[\[\[\                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          � � 6  � �@6�  ��6�   ��6�  � 7�   �@7   ��7    ��7 �������������������������������������������������������EM#_$2#####O$#?_�STTTU ##OS�����������TU #####OL9	C���������U	
**+C����������������������U	
+)*+3���������������������������������������������������������������������������������������������������������������������������������������������  � �3 ��3��  � �4 ��4�� 	 ��@3��@3��  ��������  � �3 ��3�� � �4 ��4�������������������������EMBO2#_#B#_%N# ###ST����TT��U ####)+)*+)9)C���������5)3����������������������E	3534����������������������������������������������������������������������������������������������������������������������������������������������Y���Io�օͤ���5�$ ! � ) 2   B d}�ב��ږ�Y�im-}� ( J % )  � � ��foIoKk�����j{ � � � d    � ��/�����KkY����� P J J �  I A V�fo�����I����	 � H ) d  @ 	 ��/�#k��Kk��Z[K_
 P � % �  � � V�3�Io��7��>��	 H � ) �   �  ��^_���ڥ�V�-���
 � J % J  R P +{foIo-�,n%�|��� � � R � @   #�/���em��+�֥� P J � % � ) P V�fo��Z[X�J|�S�	 � ! � # �  $ ��/��ڲ�im������
 P % I � @ ) ( V���%�����J����	 ! B I F �   ����dmY[����Kk��
 ( � � I @ � P �홽J{im����|��� B � � F    ����2������ߖ֥�  I R I   ) P Y�3{��imasJ|���$ � 	 � � �  	 d}��[��Z[����K_� 
 � R � @ ) � ��f����ڰ�J>j{H 	 	 % F � � � 2���[Vִ���-���A  � ) I @ R A eof�)�im��%��5�� 	  � F @ @ B _��������+Z[-}�  R R I � � � eo���imXܒߏߚސ  	 � #     ! _y}[��imV���Z�� � � R �  I  ��f�����,nI����! 	 	 I �   ! ����[Y[�ڬ�imZ�P  � � %  �  eof�J{Z[7����Mo� 	 � � �   � _��2�����Y�im���  I I J  � 
 eo3{%�-�������ސ � B R d   ! _��dmemKkY���Z�� 
 � � �  %  �����ޖ��R����H B ! ) d   ! 2�������Kk��imZ�A  % % �  �  �� � G@� � � � �������`��?�?���KD��@�h� ��?>�<��8��zy� � � � � � / ��������?�?�~��$ÜK�C� �h� GD~|<�<�8���v�=��� � G@� � ? ^ �������?�~��C$�9�D�� �4} �"�<|<�x����;ឿ�� � G@ ? ~ � ��}�����~���CH��KD��c� ��<�x�<�����O�^� � ��> ~ � � ������������$ÜK"�r�_ ��x|<�<�������O���  | � � y ����������C$�N�h9؆_ ��<|<z������x���  :� � � � ���������C�'҈4�؆� ��<>=������g�Oy < t� � � � ����������	�iD�lC_ �~�����������O��< x t� � � ^ �.�������ЄxɴDN؆_ �"?��O�����������x x �� � ~ / �\��0������hB<ɴ"�؆� GD����O��������=��x � t� ~ ? � �\�8�������4B<�ZD��} �����ç��������;�z��� x t| ? � � ��_�����~@��4!ɴD9c� ����O�������v���x x :> � � � �8\�����~�?@�`B<ɴ�4r�4� ����O���������x <  � � � �\����~�?�? ��4B<�ih��h� :"���Þ��������<  ��� � � � �.����?�?`�@��4�x'�"�� �h� �Ï�=���>����  G@� � � � ������?`��?@��h	�N�D�� �� ��z���8���                � � � � � � � �Ii�@
@   ��9����@� ����            ��   � � � � � � � �Ii@ 
     @�9�`�� � �A��  ��        ��   ��� � � � � � �$4@      @
��`�� � �A��� ��        @@  ���� � � � ��� � $4      
��0��� � ��� @@  ��    @@  ��@� ��� � ��� �       ��0��� � ��@�@@  ��        ��@� ��� � �@� �       ����� ���@�    �@       ��� � ��� � �@���  	     ��� �� ��� @    �@     �`� � ��� � � ���  	     ��� �� ��� @��  �    �@`��� �`� � � ���         ��� �� ��� ��  �    �@0��� �`� � ����         ��� �� ��� HH  pP    ��0��� �0� � ����           ��� �� �� �HH  pP    ����� �0� � ����           ��� �� �� �$�  8(    `P��� �� � ��p�           � �� �� �� �$� �8(�   `P�������� ��p�             � �� � � �� ��� ��   0(�r������ ��8�               � �� � � �� ��Ҁ@@   �0(�r����@� ���8�                 � � � � � � � �Ii�@
@   ��9����@� ����                 � � � � � � � �Ii@ 
     @�9�`�� � �A��            ��   � � � � � � � �$4@      @
��`�� � �A��  ��        ��   ��� � � � � � � $4      
��0��� � ��� ��        @@  ���� � � � ��� �       ��0��� � ��� @@  ��    @@  ��@� ��� � ��� �       ����� ���@�@@  ��        ��@� ��� � �@� �  	     ��� �� ���@�    �@       ��� � ��� � �@���  	     ��� �� ��� @    �@     �`� � ��� � � ���         ��� �� ��� @��  �    �@`��� �`� � � ���         ��� �� ��� ��  �    �@0��� �`� � ����           ��� �� �� � HH  pP    ��0��� �0� � ����           ��� �� �� �HH  pP    ����� �0� � ����           � �� �� �� �$�  8(    `P��� �� � ��p�             � �� � � �� �$� �8(�   `P�������� ��p�               � �� � � �� ��� ��   0(�r������ ��8�                 � � � � � � � ��Ҁ@@   �0(�r����@� ���8�Y���Io�օͤ���5�$ ! � ) 2   B d}�ב��ږ�Y�im-}� ( J % )  � � ��foIoKk�����j{ � � � d    � ��/�����KkY����� P J J �  I A V�fo�����I����	 � H ) d  @ 	 ��/�#k��Kk��Z[K_
 P � % �  � � V�3�Io��7��>��	 H � ) �   �  ��^_���ڥ�V�-���
 � J % J  R P +{foIo-�,n%�|��� � � R � @   #�/���em��+�֥� P J � % � ) P V�fo��Z[X�J|�S�	 � ! � # �  $ ��/��ڲ�im������
 P % I � @ ) ( V���%�����J����	 ! B I F �   ����dmY[����Kk��
 ( � � I @ � P �홽J{im����|��� B � � F    ����2������ߖ֥�  I R I   ) P Y�3{��imasJ|���$ � 	 � � �  	 d}��[��Z[����K_� 
 � R � @ ) � ��f����ڰ�J>j{H 	 	 % F � � � 2���[Vִ���-���A  � ) I @ R A eof�)�im��%��5�� 	  � F @ @ B _��������+Z[-}�  R R I � � � eo���imXܒߏߚސ  	 � #     ! _y}[��imV���Z�� � � R �  I  ��f�����,nI����! 	 	 I �   ! ����[Y[�ڬ�imZ�P  � � %  �  eof�J{Z[7����Mo� 	 � � �   � _��2�����Y�im���  I I J  � 
 eo3{%�-�������ސ � B R d   ! _��dmemKkY���Z�� 
 � � �  %  �����ޖ��R����H B ! ) d   ! 2�������Kk��imZ�A  % % �  �  �� � G@� � � � �������`��?�?���KD��@�h� ��?>�<��8��zy� � � � � � / ��������?�?�~��$ÜK�C� �h� GD~|<�<�8���v�=��� � G@� � ? ^ �������?�~��C$�9�D�� �4} �"�<|<�x����;ឿ�� � G@ ? ~ � ��}�����~���CH��KD��c� ��<�x�<�����O�^� � ��> ~ � � ������������$ÜK"�r�_ ��x|<�<�������O���  | � � y ����������C$�N�h9؆_ ��<|<z������x���  :� � � � ���������C�'҈4�؆� ��<>=������g�Oy < t� � � � ����������	�iD�lC_ �~�����������O��< x t� � � ^ �.�������ЄxɴDN؆_ �"?��O�����������x x �� � ~ / �\��0������hB<ɴ"�؆� GD����O��������=��x � t� ~ ? � �\�8�������4B<�ZD��} �����ç��������;�z��� x t| ? � � ��_�����~@��4!ɴD9c� ����O�������v���x x :> � � � �8\�����~�?@�`B<ɴ�4r�4� ����O���������x <  � � � �\����~�?�? ��4B<�ih��h� :"���Þ��������<  ��� � � � �.����?�?`�@��4�x'�"�� �h� �Ï�=���>����  G@� � � � ������?`��?@��h	�N�D�� �� ��z���8��������������������������������������������������������������������������������������������������������������������������������5,2?L	*+MO####O$22########O?")***+x>=>9)"	* 2
S�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������51L)+�####%$##########?%%"34445)*+)>>=<==x)9	+	+>)S����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E,%11$ht=^N#####%$##########/C��TT45)	>>==<==9))>�>)C����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5,!11$1$�=^N######/######___%$CTU	S�5)*>>x<==	9)+>>>+	3������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������45,$2%####B^######%/11$%� )S�45)>>>	
S5,345>)+ #.*+C�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������EM###B/^##B?$######?$%$11$%�O)*ST�5
	
9),S��5 #.	*+3��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E###%%?$?^#####$$�O%L�)
SE
S5***,STU #.	34���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E ##_%$_%$^%^##BB$%/�%])93U+),N#.+3�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E#%_/^2%%$??$2#%?!!"�,/#O%L9)9		,---.	
3�����������������������������������������������������������������������������TUS����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U%^%N]$%???$N####?!!"344�5?L)+C5*+)*9,-.
	

**+C����������������������������������������������������������������������������U	
S��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������EMBO^^N/111$1$#!"344��TTU$3�E)*+)*+3::5)*9)*
	+35)*+3����������������������������������������������������������������������������E	C��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5,$$_%?111$$$^%34���TU$%?LC��5)+3::5+3:U	S5)**S:5)*+3��5)+34�����������������������������������������������������������������������������US�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������TT5 !$O%$$%%$/S���U?3����5+3U	9)9	
S:45
9)**+)*+34����44������������������������������������������������������������������������������E	S�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��S45 #%%?2%$22$STU11C����E)3U	S59
99	S::5+3445)C�������������������������������������������������������������������������������������UC��������������������������������������������������������������������������������������������                   �
              s  s  s  s                �  �          s  s  s  s                                                        � � � � � � � � �                                                                                                                                                 ȡ                                                     �� ��    �    �  �  �  �o  �               !     �  �  �  �  �  �  �  �  �  �  �  �  �  �  S�����������������������������������������������������������������������������������E+C���������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                �# �# ������������44������E3���������45S���������������������������������������������������������������������������������E	+34�����������������������������������������������������������������������������������������������____��������;<=>( 
8
�





� 
(L
8Lnostefuv��������L
M
J
K
L
M
J
K
L
M
J
K
�
�
����������������H 
XY

Z[

)9 
O?I����������������L
M
J
K

N
N
K
O

J
O
�=>>������������������������jkz`��./�
)9C=D>H
XY
O?I�	�	�	�	Z
M

Z
L
[
[

____��������������������������,-lmdiBCRSDETU�	�	�	�	�	�	�	�	

�	�	�	�	�	�	�	�	�	�	_'p'p'z'q'r'y'z's'_'y's't'v'x'z'u'v'y'z'u'w'y'{'|'v'_'|'u'v'}'~'u'''_'�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	

�	�I==>�
�
�
�
r
�J�JuJtJ�J�JrJ�J==�J>=�
�
g
g
m�m��m�gJ�mʋJ=gJ�J�
j
�
z
jJ�JzJ�J�
z
�
l
 � �m
 � � � �mJzJ�JlJ�J 

m

�
�
>�
l
m
�
p
 � ��
�
mJlJpJ�J�J�J�J>�
�J>�
�
�
�
�
�
�J�J>�
�J>�
�
�J�J>

�
�
�
�
�
�
mJlJjJ�Jl
m
�
j
____J JJmJ 


q
b
c
r
s
d
e
t
u
cJbJs
rJ 

qJ
i
j
y
z
k
l
`
a
m
 
p
�


�
�

mJ�
pJlJkJaJ`J 

�
�
 

m

�
�
zJ�J�
�
>>I%J%Y%Z%f
g
v
w
m� ���



 �m���gJfJwJvJjJiJzJyJ 
n
 

o
�
x
�
�
�
�
�
�
oJ�
xJnJ 
 

�
�
�
�
J JJmJ 



�J�J�
z
O%`%_%a%4567`
a
 
n
aJ`JnJ 




 






 



1


1J

 
 
1�!
"


 JJ1� J �1J
 �

"�!�1
 � �
�
�
�
�
@APQefuv�
�
�
�













1�

1�


0

3J
 




0J
3
��V���V���==>> 



 



 



 



@APQ 



 



____



 



____ 



 



____________ 



 



 



 



 



 



 



 



 



 



 



 



 



 



���U	
STU	+#O%1$$%11$22#######################2#####%^��STTT��������5)*+3:U	
*+)+�)+)*+)+^)+ST�����������TU!�!/"I��!� ",!,)****+C������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������_____/p,_/�,y,_/�,_/_+�6�6�6�6�6�6�6��������`abcdefg


1


1J

 
 
1�!
"


 JJ1� J_/4444_/4_/ 



_/�,_/�,�,_/�,_/*,+,:,*J,K, **L,M, **+l*l*:lH
XY

Z[

)9
O?I0

3J





0J
3
4444	4
4 44�6�v�6�v�	�	�	�	�	�	�	�	(
8
�





�
(L
8L



@APQ
1�

1�


 �1J
 �

"�!�1
 � �
___P%A%B%Q%R%C%D%S%T%BeAeReQe__Pe_K%L%_'\%M%N%]%^%O%`%_%a%NeMe^e]eLeKe\e_gK%L%Q%R%LeKeGeFep�GeXeWeG%H%p%X%O%r%_%a%L
M
J
K
E%F%U%V%I%H%W%X%I%J%Y%Z%HeGeXeWeFeEeVeUeb%]%_K%^%_%b%@%a%^e[%ce`%Necebe^ebeKe__b%__be___O%Y%_%s%reNe@%[%seMe^e]e **** %!%$%%%"%#%&%'% %%%%%%%%L
KM
KK�J�J�J�JJ
KKK
�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�% ?!?#?$?"?_?%?_?____(%)%,%-%*%+%.%/%%	%%%
%%%%�J�J�Jj
�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%&?'?_?_?(?_?_?_?_+_k_+_+ 

�
�


�
�
�
�
jJ�
�
�
�
�
�
�
�
�
�
�
�
�
�
�J�
�J�����������������	�	�	�	�	�	�	�	 J�J+J�J�J�
�J�
�
 �
+
�
�
�
�
�
�
�
�
���
����
����
�
�
�
�
�
�
�
�
�J�
�J���������� ��  ****)*** **+J�J N�J�J�
�J�
�
+
�
 4447�7�6�6�__667744447_446__7_6_6�7�_6�447�4_6�__7�46�7�47�7�6�6�_____4444__6__0__4444_0_@0__@__12441�2�__4_44__44
N
N
K
O

J
O
2_4__2_4__@_____@@__7_6__@67_6_089:; 
	
K 
KKKK 
KK 
4<5B54A<5<4B5<A45<AB?9E;pqpq�0_3�0�0���������������������������������TU�SU SU #NSU #.,S������������������U+#%^%__%^N########$N#################_#__22STU	+"	
�	

�"	
��,/����"	S�������E	3U>9=	
S�5�35�,,)**+3���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L
M
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	L
M
L
M
J
K
�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	J
K
J
K
$######B!!",%##_####__###_#2###O"	**+)**+"	________�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%________�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%�%������������������������������������������������������������������������������������������������������������������������

1
 �__L
J
l
�
L
J
�	�	�����	�	L
J
L
J
L
J
L
[
 J1�0J3
 �
__M
K
m
j
M
K
�	�	�����	�	M
K
M
K
M
K
[

J J____`b�%�%�%�%�%�%__�%�%�%�%�%�% %%%%____________ac�%�%�%�%�%�%__�%�%�%�%�%�%%%	%%________***+3::5,!����!!"34534��������U)+9>3U+)**f	
S�5	,23�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U #.,.	
	
,.	?LC��U	
ST������E)+ ##$%%$%$####O>=>$__%#%#####O%?$%L)++"��,"��><D<=)+353E[\93����5C�������T�USU34:U34U	+	

)+<)SU)C����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U #.	
	

	LC�U	
S������5 #_%%?^%$N####%1$/%?_%^####?$/L	")"�=<=>� >)ST:��44�::4����TU3�����TTU>S:::U�f3U�	)
jl
 )+ST��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U #.	+3��5S�����E),_%^$####O11$/?^##$##O%L+L	L><D<=> .�����,>
3��TJT5STTTU3:TT��TU	
	


3�5<)*+=**+z|, #.
S������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E #.	C��E)C�����5),%!!!$/11$22__###?^)	L>==D<=e>e�e>e>C�US:534U	SUjl

S�U	

	+=<=	#	C�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E	C���53������U	�	
,1",11$###O^%?%??%##$%L++L=<DDD<u=u�u=u=CU	S:::TU	z|+<I<f	

B)S�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������US���E)+C�����U	
,%"M####N111^/????B?L))">>=<<D=e>e�e>eD)9		
		
9	
)*,2S���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������EMB),S��E	+C����U	�	M####%?%1122%?1L	LL>><D=<D ��d��"=D+9
=	

+9*= )ST��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5,2,S�E)3����U	
,22###_%%$/##2/1$1L+)+L>=D<<DD<,==="=D=3E
>)9)+f<	,2
S�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������EM#),S�5C���U	O####%???^/1??#####11$22)M1L"D>==DD=<D== =DD=CUjl>>+I<)+)**+=	
 C������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������EMB?LCE)S��U	M#####O%$22%????/$$#######22####%L,"=D>==<D<D< ","DD=>C5)z|>>*=9>	





#)+C�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5,2+3��5)S�5),#####/11$11$##^%?221^^$###############$)?"LD��D=<<D<=<D=DD==	+CE	>>>)+>)<S5#	*+3���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5)*+)*C���5)C�5)+)*####%^####/$##%^##O%$%############B%L"==D<�>=<=<=D��D=DD=3�E>>>>>)<9#+34����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E,)+)*C����5)S��4445)##_21$#B##_%^###O%$###O//#####B?"	+>D=D��>=DD>DDDD=>C�E)>	)+=9)***#+)+3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5,)+!^)+C����E	3�����E	+_#%##__%$####O$N###-O%?^$%^#?%?	+"��D==DD>=DD==D�D	+C�U		>>>I)****+�)*+Mh+#34:���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5,)*+"�,C����E)*+C�����E #O2###%$B/1$####O$N##/$%^_/???"">D��DDD==DD��DD���=CU*+	

9	



���<=�B)SUC���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5,"345,2)C�����53������E)#####$2%%?$$####N##^%$/^	>=����D��=D==DD��D	9	**+)9�h=f	 22)
3�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5,/"34�T�5+C������4��������5 2######???$#####%$/%"+>=�DD���==DD==>D	9	+fg
)+	9)+=�=<=#	C����TUC�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5���3TTU�SU**+"C���TUS���������U #######BN/$1^#######O%?/$$/%?^111	+"=DDDDD=D===D>DD+9)fhg)S5)*h���	*+ ##.C���E34�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������4::U�  #.	+"3���E	
S�������U	#####_%%?^1$1$#####%?^%1$?^1""==DD�D===D=D==>>D=)S5f	

S:5)=		+)+ ##.	S�������T����TT�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U ##-O-.	**+!!"3����U)S����TU	+#####O%$####_/^"	>=DD= .==>==DDD=D=>>>)9)**

S5
)�+ ##.	S������5S��U	S���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E ##--.,.	+"344���'(3���E	
+ ######$####B%N##???"	+=D== D=D==>=D=>=D>>>	C45*+)*)+9)***)*+	 ##.	S��US��4UC5)S��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������E#.			
+!!"3�����(+C���U+ #######^##B???%/12###/)+">>>>#=LM>>>>>>>>>>	                                                                                                                                                                                                                                                                �ch�����       ������������������������������������V�����������������������`������������ �@����              �                   �                                                                                                            �! E   7         O           )   �� P        o                                      ��   �         P   �    �                                           ��                                                         �    �                   �                                           ��                                                         �    �                    L�   H�   H�     , , , , , , , ,    :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �ch�����       ������������������������������������V�����������������������`������������ �@����              �                   �                                                                                                            �! E   7         O           )   �� P        o                                      ��   �         P   �    �                                           ��                                                         �    �                   �                                           ��                                                         �    �                    L�   H�   H�     , , , , , , , ,    :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    																																																																																																																																																																																																																																																																































































































































































































































































                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                c   	 Q9X       � X$         � �    A  �         @ )                                                             �U                                                                                                                             """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""################################################################################################################################################################################################################################################################$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''(((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((())))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))****************************************************************************************************************************************************************************************************************************************************************++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------................................................................................................................................................................................................................................................................////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111122222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222222223333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333333444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444444455555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555556666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666666777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777777788888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888888889999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999999::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<================================================================================================================================================================================================================================================================>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????                                                                                                                                                                                                                                                                AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA�� $ 
� � �   �  �                                                                                                                                                                                                                                            !� � �CCCCC B"� >�~CCCCCCC A&�~�  CCCCCCC A& �~�  CCCCCCC  ��   CCCCCCC �    CCCCCCC  ��   CCCCCCC   
    CCCCCCC CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIIJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLLMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPPQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaabbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbbccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffgggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggghhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiijjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssssttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttttuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuuvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyyzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{{||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~3     �  � 	�
%��    e �
!��       �!��        �!��        	P!$��     �  :$��       Y	$��     �  	�$��    �  ��� �������x����/����~������� ����~���� �����]��  �� " ,   $ �         �R�FV  C    �~��R�FV  ��R�FV     �  �R�FV  O�R�FV  xr              *      ��:���lV�1�A8�A�8�8�8�8_4Q41��E4   �5    ���E         %!"!$$$$ $(,048< �:�    �  p       �           �               ��      � ��   �          e    "#&(!( �             �� ) ��$�� �                                   �   �           � � � � �     �                              ����  
 
 � � � �                                        ��������������������������������                                ��������������������������UY| ����� ]������ �?�?�,?�<?�-?�=?�M?�]�?�͠�����`������$����?�?/��?�?������✍������?������������]�����˰˯�������� /������/?����
�����?�?�� ���H�$��K��?�
==��������K��?�
==���_y�H��}���
`�}���/��`�~�~#��N� ����K�0��<�?�/!�$����<	��$��	��@� �� ��� ?�	==���������z|�|�x`��#��=�����K�*��<�?�/��<	��$��	��@� �� ��� ?�	==���o?bhҐ?N/� ����,�<?mx��	x��_�o���$����� �����=��`�`�a���
�A�?���`��	�a���!�"h��� /���������`� ��/� � ��@�$h��� /���������a���/� ��� �@��A���Հ�Ձ����$��	��	��	��?�� �b`�A��A�?��`��4�a��5���4�4�X�4X�5:4�����54� 5/]�5� ��5�4��4�4��4��X�4X�5:4��4Հ��5Ձ�� � o�� ��������
����� �`�@�-���
��ݍ z��!���ݍ z/��0z
���0d�+	�.�/K	k�.�o����)-�(-�\����
�����o���,�\�ލ �,hҐv:,h��ph���,-��,��z�,/�h��'����������}�.��`��/���� ��,���-/�h��������w,��/��/h��
�$�Ш�/
���������:,��/��䲭ð������ /� /��N� /N� o����o���}� �|ĀoĀ?b��.��怤}���H����� ��5� ��4���X�4X�5:4�4ā˂oĬo��� � �Հ�o�4Հ�?b�4�耵����H���4� ��5� ��4���X�4X�5:4�4� ��5�!�o?bo���A�� �@�Ձ�o�H��
`�A����/H��`�A��� �A�o�4Ձ�?b�4�Ȁ�A����H���4� ��5� ��4���X�4X�5:4�4�`��5�a�o����?b� o`�a��a�o?bo�`?b�ՠ�����?b�!o�a?b�ա�����?b�@o`������|��� ��?b�(�H�4�� 5/]� �4��5� ��4�4��4�X�4X�5:4��4ՠ��5ա���A� ������o�= �/�= ��= o��	��/	���H�$��ĸo���N� /�N� /���	��/	�����(����/�Ļ�H�$��Ĺo���N� /�N� �֒�/�(����/���/���	��/	���H�$��ĺo���N� /�N� /��]�� � ���!���Հ���Ձ�o�]}�\����/(����(p�Հ����$��o}�\����?����_(�����(�Հ�/�(�����(Ձ�/�(����(�Ձ�/��]���Հ���Ձ�/��?b��	��z��o�6?b�4?b�5������ՠ�.6�4z��o��� ՠ�o�\}`��\���\�\���������� ����o�\������}��\�\`��\/������ �����o�?b���$��N� ��z��o�@�o��ň�o�����N� /N� }\(���ր�??V_�����&�Հ�� ��4���5�!��� �z4� ��u����	������&�Ձ��@��4�A��5�a���`�z4�@��uA��A��	������4����5�4�"�����Հ�Ձ�����a���`�z4�`���a�	���A�U����4����5�����6���z4�����5	�6�/�60�u������	��� ���X�4X�5:4�4ՠ��5ա����� �o�!�l�� �f�����]� ��4����6?^�����/:--�4� ���a���6��`��ݍ z6�6���8��6�ݍ z8��H��8�H��9:8�8�@���A�	���������@�-���'��������4����6?^������4��	�����������o}(�4�\�5�$��_
��6��A�`���-����0���/�� H��6����7����H��ϰ݄7����������t]��/���7����`�4 �6��7��$��� ��4�� \��5��s�H�����6H��4 �535�"5�$��C�`��6�a��7�A���@�z6�6���H�-��8��6�ݍ z8�0-�<��z6�5����=������N� N� o�(?��5	�5�6>� 66�)�4�'4	4\\��/3424\��/R4\�8\`�8��/� 8@55X�55/�6�o���=��ڶ��ڴh������d���]���_�� �_���� ���_��� �_�o���\?� �@���������� �$�������(����ħ��>�������������>���?�?�� �ڭڼھ��ĸĹĺ2�گĐ�ėĜ�ģ�������ˏ}��~����ĳ?/s_������� ��������������4��Z4�	��z����ň�?�K����(��Ą�(�ĵ�(�ĵ�Ĵ?�����_y}�\� � Հ�Ձ��!�@�A�������@��a�Հ���<o��,� -,+-,+-� �,z,�,� ��,�	��,��/��,�� �,�0��,�1_o�@��?���
��%K�/x���o�@���$���$��K���o���� N� N� N� N� N� N� N� N� N� N� � ==}\(��ր���M?�΍�,���,�?��<�d����A��Ձ���`���a�m�?f�K���o}(��<�o�1�;�0������������?���x���o�����$��K�/��� N� N� N� N� N� N� N� N� N� N� � }\(��ր�M?�κ0��?��<�?f�d����A��Ձ���`���a�o䷟(���ĵ8���8�䷀���H������/� �ĵ� �Ĵ��X��X��:�o��v����/�(��4�44�4}/K���.4�]/��o��Ȑ�}(���-��-o���8�(��Ķ�����ċ�˄ăĈć	��/0݀�����H����� ��5� ��4�4��4��X�4X�5:4�4ڇ� �o�(�
s����c�H�Ķ8���ė�
ːďĔē/0݀�����H����� ��5� ��4�4��4��X�4X�5:4�4ړ� �o���(�
s����c�H�Ķ8���ģ�˜ěĠğ	��/0݀�����H����� ��5� ��4�4��4��X�4X�5:4�4ڟ� �o��/����o#�$�H�� N� N� N� N� � ĭ��ļ��ľ���&�� N� N� N� N� ��� ĮĽ��Ŀ�������o������o���o`����ʱ`o�:�����(���`���� � ����������`�����˺ ڭį��� ��/���������`�����	���ڭ� ��o���(�����/-���,��-�-� ����>�����o���,������,����,`�,� -� >�������/����,������,:,:,�>�������/������,:,>�������/���>�������_����.��>��������4�� �,�.���-�/4��>���������,��>�����/�_�� �� ʱ ��$/�� �����o����Z������Z���/�oo�l��� ��� �M?�?�,?�<?�}����(����?���H��`���m?�� �������o� ��������x������/�����d����l���(�����/�����dߐ�䧍,?�<?8�����������}`�]���_�4�9�͏ C��	�/�I�`���:`���:�����m���(p�8����:�9�(8��9`��i:�պ4���6��X�o������z�~�ڃ�	��������z�ڏ������z�~�ڛ�	��ocQ7cccpht�� 7IM_c�1�?V�����/+�	f�����D	k	�	 -��3e		�	:	�	�	�	                 ����f���������,,,z����������y��	
�
P��tA �       !++���X����43 ������`@H0 $[jz                          �����(t� �V���� ��  �������� ݔ�~�q�L\-=Ml������        ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ������������������������������������  ��                  ���������������������������������`��� ���@���@�`�`�� �`�pUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������������������������        ����������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU H H$H$HHHHHlH�H�H�H�H�H�H�H�HINKiK�L�LaM|M��������������������                                ����������������������������������;��w�ݑ���]�`��Պ�MgY��Պ����׻��MQeܠ����y�R�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU/B/B)C�C�DzE�ESF�FfG����Ԁ�i� �������s�"��� ���� ��q���& ���� �揭�&D.�S����怞�5b5�5旼�P52��"A�&��拪q���"A�&��拪q����Z�%Ԁ�b��&�q���Sq�D&�q��SD�Dq�&�q���Sq�D&�q��SD�D��&�q���Sq�D&�q��SD�Dq�&�q���Sq�D&�q��SD��d�P� ��qD�?B�Ԁ�i� �������s�"�0�K��DK�D&DSqK��DK�&DSq�y��[�S[�5S5���bS[��.�Sb��b}S^O2��}Om��PqSDP"A#�Om��PqSDP"A#���K�!������A��A���5C��P�d� ���Mn�Mn�Mn�OqD���U�!��԰��
�����%��
毈��ˑ��
(����C��
毈���[�Ud�
�y�b��55�S[�Ud.�dx��b�bS5�K&�S��DS�q�&Dq&S��&�S��DS�q�&Dq&�q��&�S��DS�q�&Dq&S��&�S��DS�q�&Dq&S������"Ԁ������  �����C��R�Z� ���k��mS��k��nSq���K�!��Ԫ��F(=�&Cp&F(���
(Fs>��&pC&F(���҂�#[�Ud�
�y�b��55�S[�d�����
���枀bS�i�$��&�S��DS�q�&Dq&S��&�S��DS�q�&Dq&�q��&�S��DS�q�&Dq&S��&�S��DS�q�&Dq&S���P�!���0��������������D��T�d� ��"OD"OD"OD"OD��_� �P���#�����2����#����d�$�԰���#����E��V�d� ��mˌ�Smˌ�Smˌ�Smˌ�S��U� �S��#Mn#Mq&#Mn#OqD����1��S1���b����#Mn#Mq&#Mn#OqD����d�$�Ԑ�#Mn#Mq&#Mn#OqD����E��X�d� �������������������_� �V��"�q�D"�q��S����|^�b|^Sb|^�b|_�b�Sb���"�q�D"�q��S����d�$��v�"�q�D"�q��S���xF��Z�d� ��""�""�&""�""���_� �Y��mO�SmODSmO�SmP�S�DS���2\}2\�52\}2^�S����mO�SmODSmO�SmP�S�DS���d�$��P�mO�SmODSmO�SmP�S�DS���Fy���PUʝ��PUʛ��PUʝ���X����d�'����͑ss�sUU�Uss�s��͑ss�sUU�Uss�s԰�s�$����
摞�(��F
��(栏�
摞�(��F
��(栏�
摞�(��F
��(栏�
摞�(��F
��
(������
摞�(��F
��(���Z�&Ԡ�����&���&�(��&���S�(
��s�&���&�(��&���S�(
��s��
Y��P�n�%��U�
U
�U�
F
�U�
(
�U�
F
�U�
U
�U�
F
�U�
(
�U�
F
�P�n�%��U�
U
�U�
F
�U�
(
�U�
F
��Z�&�`�����������"F�������"F���Y��0�d�'��UU�UFF�F((�(FF�FUU�UFF�F((�(FF�FԪ�s�$��Pn�n��d�&�@����MM���dZ݁��	�r	P�����P�+�M12�}P���
��S��_��_�P�#�U��
7U��
U�
�U
�U
�U��
7U��
U�
�U
�U
�U����Ԁ���F�"�s��ssqs�s�U��UUSU�(�s��ssqs�s��U��UFSF�(��s��ssqs�s�U��UUSU�s͠�͑���ʠ͠�͑���ʠ��F�,���/����k���F�"���͂7�7�7͠�͠U�Uʠ�s��ss�s�s�s��ssqF�F������F�,���)8GVetVet�����Pn��Pn��Pn��Pn�F�#�S柁rQo3T̟MT6'	'6PT'�rT�k�	6r�	柁o~oT̟MT6T}�T���	�r	P�����F�"Ԁ���26��6�}n}Sq}n_5S_2MOSP5&#�l���H*9u��Wf��u��*9梱�WufWWH9��9*���u����i�����������������枑��������� ����҂�&
U&�q�&q����
�Sq�S&�s�
��F�SD(#�(#��Ԁ�p�D(
栞���p�qUF(&FU(���Ҵ����uϓϓϓϓϓϓϓ��uϓϓϓϓϓ��iԀ措s�s�%A
�摦��P������Ԁ����Җ� ���������*9��x(�(�(�(�U�U��������Ԁ���#����
s�
����
s�
�WW愄HH99汱uuHH擓WW�����
s�
����
s�
̈́�99汱uuff99**梢�������P�)���&
U&�q�&q����
�Sq�S&�s�
��F�SD(#�(#������n�@��*���qˏ�s��
���qˏ�s��
�҂��F�"#(�(Rn(͑��|����Ԁ����Җ� Ԁ��*9HWfu��x�*�@��(�99(�99(�99(�ff(WW(HH(���Ҵ�'Ԁ�s�s���WW�U�s�s���uu堓ς�ff(s�s愄��WW�U�s�s7�(�(�
�**�U�WWd���K�"�@�aa����aa���G8)��<��eV桒�({�2���<��A��F�	��K�&
U&�q���S&FUq�sUF(
��(UqUFPDs�
�qCUP����(���A�%曾�n�SF%���n��*�@�F(��&(��D��(
s�s�F(��&(��D��(
s�s҂��F�"厪�͑�%A���d[�O�����p����#�汢���汢���汢�
��(�7��汢���汢���汢�
��(�7���汢���汢���汢�
��(�7����x� ԰��ˑˑˑ��
�
����K�"�@�&S歞�D揀q�&�bSD��9f��&S歞�D揀q�&�bSD�汢��ufW��%%&S��%%&\�G8)��<��eV桒�({�2���<��A��F�	��K��s�
�D&SD��
(F
��
树sUF(U����
&F(
(�p���(#���(� �p���P�p�A�&
�S����#Ԁkmkmkmkm�F�"�@�Cnd�d���s��(.��r����������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                �������������������������������� 0  00*0  <0F0R0T0[0]0u0�0�0�0�0�0�0  �0�0�011  1-1=1  P1`1�1�1�1�1�1�1�1�122-292@2V2j2|2�2�2�2�2�2�2�2  �2
333(373G3S3a3l3t33�3�3�3�3�3  �3  �3�344'454E4  Q4_4p4~4�4�4�4�4�4�4�4�4	5555>5O5_5l5|5�5�5�5�5�5�566#626  <6D6L6[6j6v6�6�6�6�6�6�6�6�6�67$7/7<7L7]7_7n7  �7�7�7  �7�7�7�7�7888*8?8T8p8�8  �8�8�8�8�8�8�89 979N9  W9`9n9�9�9�9�9�9�9�9�9:                    ::                            ):5:@:L:W:p:�:�:            �:�:�:�:�:�:;;;;                                                %;6;D;_;|;�;�;�;�;�;�;�;�;<<,<=<G<[<�<�<  �<�<�<�<�<�< ==;=V=s=�=�=�=�=�=�=>> >.>0>B>V>k>�>�>  �>�>�>�>�> ???.?F?d?|?�?�?�?�?	@2@^@`@z@  �@�@�@�@�@�@�@�@�@�@AAA+A=ADANAPAcAeA�A�A�A�A�A�A�AB6BEBZBiB|B�B�B�B�B�B�B�B�B�B CCC9CXCgCvC�C�C�C�C�C�C  �CDD6DXDYDqD�D�D�D�D�D�D EE2EQE`EqE�E�E�E�E�E�E�E�E�EFF'F*F@FRF`FjFyF�F�F�F�F�F�F�F�F�F	G!G6GMG_GmG~G�G�G�G                                                                                                                                                ����� ��%�P��
�� �
V��� ��0��8s�Ҁ� ��W��L�
���$qU������q
�����	�`���<��/� ����,�����������,q� 
����������,b��� �������Ҍ� �� ���0��Ҵ�� ������Ҵ��� �����Ҵ���������0t������Kt����;���*�h�� ���� ��(t� �V�� ������f�� �����f���� �� ݔ�~�q�Ґ� ��  �K����Ґ�����<Ȅ���<ȁ���<Ȁ��x ��<�~��Ґ� ��  �K������Ґ�����<Ȅ��
�<ȁ���<Ȁ��x ��<�~���	����(���0�'��+���J� �����)���;� ����� ���0�o���� ����0����� ���0��o���� ����0�����
�����
��������	���� ����  ���c����<����� ��� ��P������ ���� ��H���Ҍ������  ɤ�P�
�Ҡ��  ������U���0���  ��(���U����
� ��<�x��
�
�� ����x�Ҵ����<����
+�G(����
�  ��nU��Ҁ��� �-������ �̱���������� �H�u�������������&������� ����Z����Xϲ��
�.�Xϲ��� ����� � ����� ���K� ���Ҍ� ���J�  ����� ��
���x� ��
��  ���� ��
��� ��������(�� �� 
������Ҵ��� �� ����� ����0C�� �����0C�� ��
�� �g��d�
��� ��g�� ����|�� �����0PM�� �������0PM�� �����<��� �������<���������  ���������W�H�����  ��������Ҁ��� �����
���x���� ���
��Ҵ��� ����Ҵ���� ���������	��������2���
����P��� ���%�����
��s����Є���
�����Є��x����$���x����$��$��Ҡ� ���0��d���1�<�Ҡ� �������d����i�Ҍ�	� *�0��Ҍ��*�)��'��Ҍ�	� �� ��3�@
���Ҍ����
����Ҍ��e*�0��Ҍ���������Ҍ�	�*�0ڼ�Ҍ�������� ��
��w��
�fτ��
�fτ����IXgv��������IXgv������x� ����Ҍ������Ҁ��� 
����Ҁ��� 
9����
��
��(���x��
�
<�
<��Ҁ��� x�y�M��`P� ��(� ����T�������T����Ҵ��������
��F� ��������
�����T��.���8�T�� ��<� |����
���<� |����Ҥ�	��$� TF��
��<d:���� 9���� H����� ��$@P������ ��$@P����
�� �����(tY������
��� ��d��H,����.��<�
����T��Ҵ��
��r������� ��M����
�� �������0���
��0�
�Ҡ� �� ��*�d�Ҵ��� ��9�d������  c��7��L ��7����������L �����
���t�  �z���Ҁ��� ���S�Ҁ��� �����D��Ҁ��� ���(K�Ҁ��� �����(K�Ҁ��e����@�������4[�,��
�0�������
���4[�,��
�0���������� q�&�`�� q������ 	q�&�`�� q�����(����g���x����
����P���
�Ҡ���*�	�������P��A
Ҡ��*�����Ҁ� ������ ���������Ҁ� ���� ��������������
�
��0�������
�
��0�����:��(�� ����7���������
�
��0����������������������������������������e�������������8����#���������e�������������8����#�Ҁ����;��
��(o� �Q�������(o� �Q�����0֐��.�������0�֐��.����vϔ���vϔ�� �����<��
��  �֐M�����
��  � �������`���0�D��`��@��A����
���`���0�D��`���@�A�������˓̱��������H�u��������0d������|� �� �������0<� �� ��������,� ������������ ����� 45���������$
� 
������	��$
� 	����(� ������� ��	��|�������<������� ���  ���������  �����3��Ҍ���`�7�����������Ҩ���3���`���`�s�������Ҡ����D�	��  ����  \�	�j���  \�	�j������(~�x���:�i����(~�x���4�i���� ��
��0�
���
������� ��
��0�
���
���<� � �<q��<q��<q��<q���<� � ���<q��<q��<q��<q�����  ��0`z������  ����0`z��������� ����
�
��������������F
������`"�ӌ � �+���� �`"���ӌ � �������,	���@P<��	���<��Ҵ����b�	��Ҵ���X�	��� �	���;��,�;�,������P�0
�	�����������T�0
�	�������5���7��x�	��,�;�,������5���7��x�	�� �,�;�,������
�T
��0`5�`?�2�Ҵ��9�����ϓ����2� I�`������6�`���� � ��m���� � ����m����������*���������(*����
��Xϲ���Xϲ�����gh��	����Xϲ���Xϲ���������� ����	�������
��  ������H������$����$��������$<����$�����
���������������������������
������*��*����*�*�����0�P�������0�O���P�����`�������0���P�������0�m���P�����`��������0������3���Ҍ���� ���;����� ��$�������� ������������
��h������(������Ҥ����	�@�Ҥ���	�@����
�����I�`�o���
��d6�����
��9	������
�<G�PV������
�<G�PV��x�e���x����� ��� ��d �������� ��������	���E��������� ��� ��`0�����`������҂���� �t)t�t��� ��� �����
��0<��0������� ���В���
��0<��0�����Ҡ��� ���@F� ��������Ҡ��� ����@	�F�� � ������������**��Ҵ����������Ҵ������ ���� �������D� ��𸥵�����
���
�	�����H������
���
�	�����H������
���
�	�����H��������  �K�������� (� ������Ҡ��� �����֐������� ���N������ �N����
�� ���0���0�	����0���	�
� �����0���0�	����0����� �0P�
5������ �0���������  ����"�֤���������  ���"�֤����Ҍ� �0P�
�
6����Ҍ� �0��
�������Ҡ� �� ��0��@��k�Ҡ���� ��(8p�Ҍ���W��O�Ҍ�����W��O�Ҍ� ��  ��H�� �����!uu�l�Ҍ� ���  ��H�� �����uu�l��Ҍ��� ���e�����������	�
���� �����	
��� �����	
��� �������	�
���� �Ҡ�
�+� ���.��2W���Ҡ�� ����6��8W��������	��Ҡ��� ���9	����������������������
�������*��*���*��Ҡ�� �����Ҡ��� ����
���������� ��������� ���������� ��������� ��Ҩ����Ҩ�������Ҁ�����`����Ҁ�	������`����Ҁ�����`����Ҁ�	������`������҂��� �*9HWfu�����҂���� ɠΡ�uW�k����  ���u���������1�����ȭ��Ҡ������	���x�� �����x��� ������Ҡ���x �	H�����Ҍ���Ӏ �HWu������d�������=�����
�
����0�D��H#2�,������
�
������0�D��H$2�,�����x��~� �� ��2��|��x���B��� ���@�Ҩ���� �fu���$���Ҩ��� �fu�����Ҍ� �� ��2�Ҍ���� ���P�Ҵ������  ��E�(D��(���Ҵ������  ��E�(D��(����x���<�0�Ȕ���� ��0�Ȕ����x���<��0����X���� ���0����X������        �4DDT3TDC�|������̋��������        �l������̊�������܋��������        ��̼����܊���ͼ��̋��������        zS2"DDBz�����z������ z?##2"$zD2"DDB{����ܼ        ��!��$/�#���� �B��!��$/�#���� �B        �l�������        ��̼�����        �.!�/�B��@�e����G�S�4���.��"�=���ڰ �cΪ2�/�S��3��/�� ���c��o��?��ER� #�3�L ������O��!.�1֪=�<��=�1 ����4Ы�Ͷ� �R��P���PҺ���!��C��EQ�$�!�\֪,��R>��_���#�P�?����<�uʶ����!�� �� d�4��c�D��3�.�0Ϫ�Q�/?��=�A� ��#�3����#��,��S��C`���B�0����P1��A��Q��?�� 1��Q�$�R���o�G!�_��3�3�Һ.��ܶ�1��1��MѦ43B_��˺�����0"���-�A#���`�%@��T��0%?��0�A0�?�C����b��� �[���3/ߪ �3�� ͖��1��l����� ����� ��<�?�0�B���^�C�4���� �3Cͺ ����@�@�^���0���!���.��Q��@�d� �        ���C��A��%�R�!��4�2"�1%0z�T��5_�z/�62���!��C���A�� ����� ��� ����!�z�#��1�V���C��!���1��B�z�O�4��3!��# �$/ߊ#"�B!z�W<�s��� $.�#�  ��P�CD.�51ۊ3��0�����Dz��/�6N��4/���"� ��B�����Ί��!��2��� ����� �������!�����?����C���#1���        ���`�"��!3�����u�1�B��D� �S���`���1����=��A��K�A�;�0� �.�?�0������#��=�/�/�� �-�2�A��B��4����� ��3� $�P��D1�����O��]�\�]�L��c�A�?��2�K���S��4�� �"�/�C� �#�/�@�0�� �q�"��!3��        �Sc�6>�#�Z��5�3�Ơ��L�E��o�.S����".���<3��'K�"���k�=!+��®2+6�_�¿<���s7�-�b�Cf��� ���3�Kߙ�@4�`���&�_�E�Bc�6-�4�Y��5�3�        �  �!ۚ�2!��=��O��Fb����C��/��S��"��"�2?�! �  ��@�3����0�1��1��E��a��F5O���S�����S��@�����#/ϚV��  � 4�1 ����A��!���"�$ ��ߊ���f � ��C���"��D@�/ ɚ��C��@ ���5�BT��龊 ��Ec� ��0ۿ-����t !�������c$������!�6d.�C�����eS�B�������Gc�%!������5��C������֚a  !�����e!"#�1�����e!!"2��͊�ڽ#d2#�!���˾#�4A2�����D2�"�����C"B���ܾ22#�2����!�#" $A�������2!4�1�������2 D"������2$#�B �����1 #32��۽ #D�1 ��� �!#C"����$D�����z�Gtf0 ����24�B����D2���� �3�2!"�����4B" ����� C�"!#/�����3"#������3�!2����z��5US%w@������#"�11��ܾ��2F=��˼�$S��/�e?���� �%B� ��� �s 0�ܺЊ�4#"1����� �C3$����5C�C�ͺ��2$B$?�컊�  �Cd�#ۻ���3!4D@�뼊��!DC�1 ܻ���DC"�ʊ��! "D3�1������4D!켊��!!4T�"���� �523�̊��� 34�2 �ۼ�!��"33D�����  24�C!����!E2"ۊ��S�4Aۻ�� � #3E2ˊ����"$�T2˫�� ��DD2ʊ��� 3�ED���� � DDS܊�����USܻ�� �  FC ܊���    #�DE0�̼��� �ET1슼��� �Ee!�˽����DUA������  ��FSB���� ��4VB������ ��4fB�������5eC����  ��5UDݼ���  ��5UD����� ���DEd.�����  ��#VT ���������#VT �������#ET1����� ���FT!�����  ��Ed1���� ���ED3��ߊ� ���EC3���� �����DDB��� ���D4D����  �ߊ$TC ���� ���$TDzNܩ� �̊�#EC!��ފ����#ESzR����뼊�DT!�ފ ����DEzc�����ˊ�EDC�ފ� ���4Ezu�����ڊ�4T2�ފ� ����4E�R��� ����#UC�݊������$T�C���� ���"ES �݊� ���T�C ������ED�ފ� ����D�D1��� �����5D!݊�����4�T!�������4D2�����4�T1�������4DA���  ��� $�D2 ��� ����#T2�������$�D2��� �����#DC �z�� �̫�F�DB�� �����#D2!�z�� �ʛ�5�C3!��  �����4C�z�� �ܩ�$zguQ�� ����#C! z�� ۪�zWuC/�� z���WfCz��ڻ��zEfS��z̹��EVTz��뫬�z5fS!��z캬�4Vc1z���ʛ�z%UE1� z컺�3Ve0z� �˚�z#VdA� z�ʪ�Vd1z   ���zWc2 z�˺�Ee1z  �۫�z�ET!!�zܺ�5T2z �ʼz�ED2z�컼�5D3z�!�z�#D2z �˫�#D2z���z�D"! "z �ʼ�42z!�˼z�32!!!z!���D"z!!1��z�#2!#z!�ۻ�#3z!!ܻz��2#!"z!���2#z1 2"�z��"3!z2���#z1#!�z��#! "z����2z!3!��z��2"z"!����#z!3��z��2z3����"j14UA�z��"�#z!1�ܾ!j"4TC�z��!�z"1����j23TDA�z��� �z"# ����j�#DER�z���!z21���j" !$fS�z���  z2"���jfSz���   jDFT���j Wej���  �jVu.ɛ��z  �33/j�����jEf1ڼ��j� �Fu0jܼ���" j�6v0����z� ��$Cj�����"�j�FfQ����j���6fAZ�����?�j�$fQ����j���%f1Z�ʚ�3�j�&f2����j���%f2j�ܽ��j�eC��j���UBj۾��j�VB"��j���TDj!����j�E4B�j���DDjB ���/�j�5B%?��j�$ ��TjC��$0�j��C6S�j�D���%DjE1���2 �j�� %e2�j�"���"3jES��2�j� 3ES�j�1 ���!jES��$/�j�  ET��j�4���z$1����j�� VC�j�0����jVc��#!j���Wc�Z�#S����jUU-��?�j���Gc �j�"����jFT ��!j����VU/�j��ܼ�j6T!���jۭ�Fd �j�̼�j6u��!j��%d j� !ۻ�j4C3��"jܩ�DD!j��"��j#DA�jR���%T"j�#0ۻ�jC"0�� $j0۪�#2#!j��#Aۼ�j$3� 3j1���31"j��#2���Z�vFe�Fj1����#3Cj��$2���j�"$4��$j2����"Cj��#2��Z��Fv ��Fj1�����#3j/�#2���Z��Vt?��FZt�����6fj ��42��j��D ��5j2�̽�3j1��51���j��30�4j1 ����4j �31��j��3!"j"���3Z@�$UB�j��3  2j �ܼ2ZQCC��j���2! "j"!�ʽ�3Z@42"jˬ�3 �/j!"��"Z/C!#D+j��" !z ��j�!�Cjʽ�" "jD.���!j  !�$Uj�� "/j�Uʮ�j/�3�$e/j�����" j�%fʬ��z�3j˜��1j�%v/ɬ��j�"��5VOjʭ�� 1�j�$e@����j�!��4w>j�����"�z�D�� �z��Cj����#"�j�gB����j  ��5fAj�����$?�j�&f1����z���#Cj����41�j�%fB����j�2��$Uaj�����# �j�e2����j�/��VAj����#/�j�f1  ��j�$ܾU2j���j�UB��j�" ��D2j/����j�U22��j���C4jB���  �j�E42��j�"/��4Dj3!���?�j�4B$1��j�3 ��C#jC!��3/�j��"FC!��j�3���$DjE1���1 �j��$U2�j�#���"#jES��#�j��"FS�j�0���!jEC���#/�j��ES��j�4 ��� "z$1�� j�� eC�j� ���jVc��2!j���Wb�Z�2S���jVT�� j���6t/�j�����jWS!��"j����VE �j��ݻ�jEU �� jڽ�Fd0�j��/ۼ�j6e��jܻ�5T!j� ! ۫�k4S2 ��2        j̮Uk��SKj��d^��z20�C^��zR��c
z�Q�.�1ve��3%1�z��21�v� �$ ۽%���#���R�D=�"/���!��#N� �  �@��z>�#�1�z#Q�$�z���!�/�!�����3^����a������!�Ma���� %���2�0��$����#�"C*�Q��B�� �0�!/��2���# ��C��"�$`���$ͦb���R��2�� ��C0���3?�1ۊ�2� ��$�##�3���2�_���c��2 ��B��S�2��d�a�3M ���4ϳ#��� /"1��3���� ���"O���  ����VN���#S����# �b���S>���C����N����A���TK�%�3���g/����D�� ���1�#�� ��� � �"0�� ��>�b�����+�/��=�Q����A���"�3�#;�!#F��0�/�B������?�C.��?��"��b����0��"�A���dߊo�C�5BL�� �S�"��?��!���D-�����#���d���1��A���E�� �2Q�ߟ��1#/�� �0���#-����`�Q����5/����0���VS �� ԊR�D���FP����V
�/����#!������PP������4��/���C?��5�"�N��12���3>����5�#-�� .���B��4 ����S>��-� 4��#�$/�ߚ#0���5�/�0��/ �,��# ��N���2 �Κ�D �?ۚ�#-��D� � ���C���$1ܚ ��0#���32��@���3B��!�3!��/���3,��$2��"�%2/���#A��?���1.��C�2͚E ̽"C���.��R�O��#��4��4O�� E���!�!� #��%>��1���&Mъ���#�rښ��1�N���2���%Q���  !��%
�.�S�]�v����D����c�����$0�d����v��@�D���1��d�����2�#����fO݊�2
�6?ʚ�d���>�5�-�ޚ2���#0���U>���3�3����C�"� �P���50��.��1��D��!��C����C�0��#�D�� E?�A���r���2��!�"��#� _ޚ�"��4��� #��!���O�".��C��"���$-���C!���R��#�� �B����4�� ��32�WQ���B��#� ��S��� ����T��3њ?� �̚C���!� �!��r� �C�?�"� �b�њB�#�E���4�PΚ��D���2�3���b��R��Q��3?���r��1���C�ߚD��R��%�0 ��E ���3�!��A��C�C���EO��ߚT1ܰA�#���S��#f��"�/ � ��2
�4���3���0���"#�2�ʪ0��"!��B/���"۱S@���0� ���C�/܆�EeTVM�� �! ��A����6��B1��1 �����@$5.۪��A� ��#<�1��3�N���"1��2/��$T����$.�3���S����43���B��!��2?��0��F>ݚ��3�%R.���CB��#�� �!�Ϛe@���4��F3 ��51��%�1�� ��&P���1�@���T1��D=��"��5R���S��&c�vO��d@�Ҋ��U���Q���b����A��# �޾T��3����A�͚C�T�����eO����1���!�0���b��S��51�њ0!���C���!�0���T�� 3���A�� �њR�� ���B��B�!��/�C�� ����f��=� �t�Uٚ��@�!��� ���3�#� D�� �T����a�/��$$��B��"���2���3�����5"�" ��4B�ϖ.�˰B����B ��"��&�TR��M���@��$��,�# ��f �e��!��o���"?�� �4�W��5�#�Q���2���#���A��C�Ӛ��0� ��7��d��B��0���/�&�ϊ0"����%T��P�T���2  �?�����Ú �#�1���C�݊U��� �� �4 ���A�"� >��R��=�&
�@]��&.�4�� .��V���0��1���D/���BO��!!.���A�� ���R� .���"��� ��C����B��Q����"/�0���Q�"�ѪB�����!����/ܚU�R�3���U���!���P��5�Ъ!��B��5>,��5P�� ��B��"��3��C3���A1��/����@��$��D+���#?��" ���4����"B��@���3Uڡ�U1���d����1��� /��@��3�� ��5�3.�ߊTq��2�#���0��B���/����0�� "2�2��$��  ��V,�� B�-��B�ݚ%@��d`ͬ�S�� ��� -�C����#�!��1�������UM���A��3N��""��"1���2�" �Ъ  �  � ���?�����#0��?�3^��"!��3 ���.Aܬ7� �/����#��&�-��1�&?
��"0� ��#?��4P���D���W1̛6 ۊ7�A�_ڪ  ��T���� ���CN�� �2��#@���R � �#0��� ���A����C���0�� � ?�1�E���3��e���##Q���A  A����c,�#ޚ!/�.�DC���$��#�"��F��2,�C� �.��1����$����D\�.�c���2��C��6_�>���F?���"���Q����1�DN�����A�1��b��1���" "��C4!��� �����1ܖ�B��"�"�##2ۚ�5���D�A���#�""�#0��d ����S�0��VI�AE�� ��$����gۚ�0 ��Ϛ1�$e��B� ��D?��0��R;�E!�F��1���� 0��E-�42��!��"3͚"7��"R�=�"D.�D1��/�$њT<��EN�̪!�����R�� �!����$�.���U��� �5B��!�3�C���$1����FI���,�C�� 2��b"���3>��0���GN�� ��4B�$<��g!�@��#=��Ua���� ����B! ݪ"���#��$"��!�! /��R��C?#0��23횽�T/� ��$R���� �0���3?���#���� �A���2��B���D ��КTc��B���f���DL���2��C!���3���.�S/ ���@����1��3�C�A�� #� D��Q�� ��C���3.�ޚB!�d�Қ2�����VP���6!��=��$�.��#2!���1��q�� �.�"� �%b�E�� �d���  }�� /��2���DC��@� �C���#�!��4��!���R�  ����TM�Ū!!��3@�Ѫ"��"�� ���$���3��"��0��3��$���$O��1��#1��2�� @�ܪ!���@���R0��c.���2�њcܳs�޼�S��#��T��"���$��4����B��SQ��!3ޚ�1� �EB���#0���4�0��4C���4/��1�@���!��1���4@�24��% ����!�"ۚ�v��#��"/��@����c��! ��"?��@ �0����B����2�!���A��P�!��o���U24����E!�"2�ݽ�B��@��"O���!""��2B��� ���"��P��/@͚!��""˚�#$�O������4��O���B��4 �N�1���4`���"%b��.�� B����31�?�#����!��"B�١.� �@��## ��#-��5P�3��/��1�.��$�A����� ���#B͚ $0�1�1���4R�?��  �5�AN��%_�3��$�� %S��� � ��$1���1�"M��2���!����1���0��0� d���?��۪1 ��O��!e���0͚��C �Q��2��$4-�����_���!���2��b޽43 ͚��A��К$.�!�� "�/,�C��1!����"A����W.�.����U���B�Ϊ ��#?����� D��U-��""� ��D ڪ�% �����E,�6 ��#0���D� �30���Q���6.��3A���E �����$�C��C����_�$!���&_���5���21���A����a�C1� �0� �-��W���T���Q��5��4P�����К22��S��>�S�V?ښ�%1�� �� �Ҋ4/�.�@�R���@�Қ0 ��!��?��!  ߚ�A��"� ��S����R�@���� ��Q��#/��4���1�����"1����R  �4/ ��#���3���A���"����S  �� ���%M�̪B�! ߚA���d���#?��&�/���E�C����!����CDC4C��$?���S�/�2��� �"��D� � ��!��̡f?�T�ߊ��#T�E�d�'0��R���%2�����A���S��$O��ߚ!/���A���.�"�� �#���4/ˊ .��t�1���2�?���F���5.���B����U<���_��2���S ��.��#6����d.�^���" �3���� ���T,��0�>�"����b���.���!��S�� �����C�� �!/�B��%B� � ����2���/�P��4��5@��_��5��<ҊC�$����� !�4��U�/�0��<���v���!���2����F��A��#� �%��-���2��/�$
�D.ޚA��>���5.� � ��C�;�e괚4-�2��"� ��>� ���d�
��1�"�B��  �� 3�0��� �S����C�TC��2��1���$ ����3���QΊu-��a��. ��30��2����`�4��0�"���5� ���$0�����1�3�� 1>�T���E.�!���%0����B�5��#!�! ���E Κ��E? ݊�E1��r� ����D?�/��V�  ���1 �0�#1 ���3"�N���6@��� �R��A������20��1��G!���C���1�/�̚�1�@ۯ�F@��T��0�>��.��0��"��F"��E�/��%� ��@���0�6@���! 5-��2/�3��O���0�� ��E/� �3.��3���2�A�����$1͊�? U� ��1��@��S�/��F� ���"���RP�ҚA�? ���%�A��N� 4#E<�a� ,�`����N��0���"�D��3 �����-T��@���@���U�c�D)��]��C��D��2�3�F���� ���S��R�����"�E���/.�!� �?��p��d����Q�5&:��!-��� ޚ���3���=�/�!#�,�.�0�0ݚ�?�� ��/�T� �0��1$��R��!��0���1��-�dЊ_�3�%DK���S�"��N��!����U�!�"� ��e���1��@͚�F�  ���"a��A ����� ���#.���#��P�R����E���%��~�US��!�ԊR�B��GP����V�/����4 �����`�P���" �%�����C0�!%A���S�����3C���3/����4�#�� -�        @�� L�."�  ����� � � O���QM�#� B� =���O2�P�Z   ��#$ZE��A��Z3�"�/Z��A�Z<���N��j�4��@�=z�#.��4j+�0��S�j�B�4 �&z.�$N�$/�z � !�%/z��b��_�2v��C��E?��>�"���?�"��$�.���v�/O�4�%��!��0��v��M� ��D�R��z0��9��R��1��� �4�.��P�N�.�Bz��2���3��@�B�����1��!�2���a�<�"� �@��$-��U��B�R���D��f���3�D��0�z�e��"��2z�"�-��.�"/�$-��2��"�"��"2�?͊#�%,�6,��4�R�$�� �.Κ?�5�  ��4�1 ��A� �0ݚ?�0�.��C��!���a��2�Q̚ ��2��!���5�Q�Ԛ1��!��!���b��!��A��!�� �$�dڊR��#���$>��F�"C���2�1��P�1�e��C��$/����@���C���MŊ_��O�0���O�b��ՊO�$��3��DEΊ �!��  �$0z�������D��C���1����$?�� $1"�����6��!�@�B�bۊ��6M�?�� �4���@݊$��B��O��40�����U���2� Q�����1���r���&S����� ��!��%�b����1�����B���GQ� ��ъ1���C� C� ����!.��2 ��G_�� ��"/�����4/���V?����Sz�
���R����U1 �����A���5�>��$C�����!�$�ЊC�S��3��#���.�D/��e?���B��1��3/�B���U!"������3�� �f������a�.̊�#�ezq����C���#! ��S���Њ2���T�� �&Q� ���p� �ҊA��3T�� �� Aۊ���3�"2���#-��$ ���4!�����!���C� ��C���A ���2!��C1z����E2.���A��&a����?�� /���U!�Ί@������&b �����A�ߊ�!��$S������S���2�Њ61��A��4��2��&s�݊�0���� ��C����EO��� �!��V� ����@���?̊e���� 1��  �C��C2�ߊ�$-���!�C��C""����# �z��T1���U �����C��$/�� 5B����0����!�4Sފ���"͊�"!��V0z �����d���3ߊES����zE1�˼�t�� U ��z��Eʮ�" ��!R����� �#���"�Dzs������5zO���3! ̊4C�����2��3��C3���� �! �ϊ#�/�7b�z����6-����! ��e���  �0�� ��D2����z�F0��2�"�D"�����͊���5Cz������3!zʽd�zFe1�����z40���cz��EfQ�ܭz �3��ފ#!��2"z���2�z�E=�fze>�����$z@���%R���#D��� z�$@���d�� #C��z���4!��͊�3��S z�����1�z���UA���43��������!��41�������!�"�42�z���30�̊�2��42z0�����%Ozܻ�$T/��#3!���� z�B��d0���#S ��z�"!˽�"!�E1�z����1.���#0��Ezc����"!z۬�4C݊�EA����z�%/ʭ�2D��5R���������$Cz����!܊��"���D/���� zAۼ�S!��S����z�"���E� �T!�z����C�˽�"�T z����3z���#D��E0���� z/ʽ"D/���C2���z  !٭�!� ��EB�z��� �̊�"��$Sj�˚�"$Ozۼ�E ��D ����z ���E ��$3!���z��!���!�T z����"!���DzP�����3z��!#C�41 ���z3���#3z �Ve��z��!���!��4Bz����"ڊ���3�B����zܬ�#2!�� C ����z�#!ˬ�C� �C ��z��#/��z3""�6f0z�����#1�z˾31��D �����z��C1z�$gR���z�"1����C� �C! �z���3˭��$2z����"zܼ�52��3B���z4ۼ�32� C���z�# ۫�3�!  �#3z���3/��z�C�Guz0��۾�4/z���1�D �����z"2��D � C! ��z�3���# ��41z����#C���"�4zb��˰4!z ʽ�D1���$C����zRݺ�T2� �4B�z��3��"� E/z�����30�z��$B���C!���zR��%S���D0���z�"3��$B� �D1�z���3"���1�C1z����3.z���E1���42 ����z#���3D?z��fe �ۼ��!���"��$C�����!�Ί�"��$3z0��ܼ�3!z���$D��D ������2���2��4! ��z��3���2�41 z����B�z��V@��gzS ����#Bz��FQ��$3����z�D���FR���34/��z��20ʫъ#"�#Bz�����3 ���1 �#�D/�����z0���6S���T0��ߊ "��3���D1��z��#1��Ί3?��42z����Dz���FR���E1����z2.���UC���U"���z�1ٛ�U�!��4C�z�˾4/����#!��$Cz/���2z��$v��#D ��� �!��""���$B ��z�1��#�"!��$C1�z�ܬ�#2����#!���Uz0����� z��6a��E1����z�4���ER��D"��z��#.���"��5Rz����?ʊ��#1 ��4zu/����!z"��$U?܊�4C����z4?۬�#F� ��S��z̿"!��"!��Sz�����1�z��TB���T����zA���#C2-��C"����z�!��U�!�D! �z���Bʽ��"!�E0j����Vzʽ�$T��D1���� z/ˬ�#D/���42 ���z�  ʼ�2���62�z���ܼ��! �3Sj�˫�Rzڬ�"D0���D/����z���D!��#C ���z��# ����!�D z����"����Cz@�����3z��33�D0 ����z�$���"Cz �gd��z��"˽���DAz����"ڊ���3�B���� z���#3��$B����z" ۻ�4� �$C�z��" ��z#2�&f@z�����#!�z˽C!�$�D ���z��32z�%gR����z�""����C��C! �z���!#.ʝ�"�51z����"z̼�#B �3B����zD˽�#2�#3���{�3��3        �   ���#jaA�T�	�� �� ����E?���d�D  ��%D ۭ ����/��!�#���B���S�B��~� �� ����� �@ъ A/� �/##����4�.�ފ�����ЊR!���`������.��2�0��.��� ��zF% �$�O�@�! /�.z!��������0zT���Ov�����z��?����z������Sz".��B1z�?C�#z�/�!������� z@1� Az�a !�z/"����z������ zQ0��zC !�!�j-� ܭ�z������#zA�z0$  �j��^�ݻ�z�����"zT2��! z!0j�A����z����� 3zD �  !j$D? #.j��12����z�����"jFR��4Bj#!E1�j������z���� "jcA��0#3j%B#"/j�!����jʪ����VjS"��!�#0jB#/@j"1����j�˫���CUjB��#"21j�23!P�Z $ܪ��j����3$jB�j$B##!2j#�����jʼڮ� 5SZ!��d25jT!#C3 j21�����z�����2j#-�� #jDC%!$!j�����jɫ����2EjO���3#jBC 4!j1 ����j������DDj@��22jS3!!#2j �����j�����E2j��%jT#"#2 j2/�����j�����5Rj/���2!%f�2""ET2j2�����j������5Rj���25g�"""UT2        3#��b� �j     �lZ�� �N#J�AP�C4EZ�A�/ V� AZ ��2V����Z��?���J���
�V��!ZS��! >Z�1��O$��5=�e�3�g�^4� ���в �����N�������� �M���1�q�
7���.�2�*�3%�!���̶"�Z�-���!� � �/��@�� ����=���l��9���C<�4�@��@�0�#���D�O�Ҷ? /��3�E�4+���?�-���#�l�+�������/�.�/!�!�>�. �"C �31�2"C�?�!�/B���4����>��������OݾЦ����� ������!��#���!��1�/��"��� �Q��.#��O�>O��l�Ac�P��p"�"�O������<�� ��� �C��-2� 0��!�-!�=�/�2��$��?�"�0 5���#���0�����!�� ����2����!�����@��,�������� ��������Q�ܲRN�!���E5�"� ����B��.��>���2��M �]0��T?�D�>�T�S�2�\�o�.�c�L'�6^��U�.O��/���������#�P� ޖ������ښT�@��L�� ��
��/���Ԇ��>S���?�!�B������!�R�������O���"" �0�"�!�M5,W�%�b2�]�1�@��>�,3"1 � -�����1�"�.���"����-���� �<���� ��BݱL���/�3�� ����/f�>ҖA���� �e� ���=$��?�����1�&n��-�d��# !�`�E�4L��d�@"!�2ݚT� �-��M��?���O�!���������@�-��/��/���҆�;�,���� .���<�O�  !�4���@��.���  B��=Ζ���@�Ֆ�����N���@�>�4��U�EQ�@"�@�%�#]�$/���0�! �����U�������M��A�?!����.���."�?���d�?��b���Q���3�"��3a�K�ݖ!�7 �������#>н�_������Q��@�?#���4�2�0 !��@m�3��n�21^��2�@�4�P�>��0 ����� ��� .�
0#��*��%�$�������
����"R���?��� ��S!��0�D�C3"A�o�`��D � ��0�t�K����/�1>��"���C��?�S���5��P�<�<�\��C�R%��S�@�A͖��$��"���2���U���� � /���R�� �<���.����-����/������!���?��.��A403�E�,����5�0�-��O� �ߖ ��0�� �!#Ҫ� �N�?$E/і2D�T "/���>��>�4�%�!���?���2����ƖN���� P������"������A$����4��.��D�/æA�""�,��        �=��!��0��R���#���2�*Ԋ�$��3�>�"��a�@���N�  ���_��ц?�4�b�1�L������O;��!M��܆��6�$$B�k�T����̆��.�3$,��� �?ߊ��C� �� ��L�,����0�A�.��!܊0�#�R��#0�0�����b�$M�N�#�1�������?"��� �@���"�O�s���?�,՚"�����@�/� �����12�O�.�ޖ����>D��1�o��"������C�/�  �Q�@���� ��#��# ,��<��"��/��0����-%͊B�M�/�0�� �,��2�!��O�N�E�_�{�M��"�! ��S�"�����$�B�.�O���0�^�b��G)�Q���?�R�4�� �>�0�"�������D��5N��m�����L�� �M��w��!�>�.��Q�B�.��-�����,� ��B�/�/��@�!���3�2�@��z� 	#Њ�2���Fe0>��������0�
 ���?��A���/�?��$݊&��n����0�0v1�+"#CDz�B��� �>��1��O�P�-���P� ��.��ܖ�������!�D�2�@��>�a�0/�O.��Ɋ  �3�!z�?���".���>U�U�O��@�O����r��� �? �D��!5/%�n� ������� ��D��/O�����/�=��?�4�����"��'���?���O��]��d�-�n��]���3N�@����#��D�=�@�. ��2��MÚ,� .��!�B�Q��0��"C�  ����#�Q� �B 5!�
����S�QE2�D�P��� ��>��p4! ��͚/�2�0�l����0��{�M��#�"D!"!���#��->��"����-��!�+�z.��s�M�Q�#�_�p�������"�>���A����   �-�ޚ@�1�#��D"4D0�N���  "� �5*���=��o�1��^К��!�/��/��@� ��>�����3�?�� ��."�#0���?���!��?�����@���-��*�N�� ��� �M������ ��� !�"�Aޚ$��,���J�6��"���#�"�1�^��k��#��b�#O���� �3��"����#��1�>��=�� �����M����0�AV151�3� �9����#���1�������^� ��0�2��A���&�"�?���&:��S�� �!O�!�cA� ��Ж����/4��D !�����/�2�"� �O�A��?��V���[��1�?���4�.��p��02��0�p�3��!��B���������5�m�!��@ϊO�B���#��3� Ϛ0�< ��"�\��1���<��$��"�/Ҧ�����2��B!3���̻�ܽ"���.�"�M���0�2�|� �"���!�1�/�� �&����.���O�L@�<��3�2���_�B�/��3���:��� �"�!���� ��%UUVfW]њ � �A�0���>���d��,�,Ӫ �  ������%�$��1�!�R� ��]� .�c��L�N�� ��=�O��0�*��0���-�� ���� �� ��`�_�\O��.��.�.��$�!���� ���/���Oߊ�!��T���!�n�?К�+��.�.�'�-��A�/���=�.�/њ����� !��]њ���/��B3,��A������,�oߚ�
/��4�"�!���! �����2�/�R����>� D�#!��"�.��2o�!�/3���1��3�.�S������D���@�N�`К�.����U�^�&��O����O�O�2�M��˼��D�4�"�z�-ܽU��?�>�6��-%���u��O�b�V���-��?���!�<��s��1�� ��2�>��C�#
���2� �����!�1��$���"������2�"�O��<� �"��<�2�B���� �+��0�C�,�� �R� ���2���^�+��0͚�,%��������#2T"��$�2�"�l��/� �0��2/�
����"�"�3�Q��"�/�����  ��C̊ .��2��]�U�P��#�������#�@�C슱R� �!��C��>����������K#�c�<���u��_Ú�1�.��V
�/�O��"�0��"����$@��$4��V�@�M�-���� A�D�<�N��?њ�M�4�"��c�! ����"�/�Qߚ �n��N��_��?�.�.���������C���9�6��2�.�!z��O�j�1���"� �b��)"����5�1�3ъ[�k��� ��E�Іb�T�!�έ�y�-�&��_�0� ���e�C�@ӖB�"�1��ϊz�-6�P�>�&�P�������!�C�/��݊Q��!.�Cߚ!�?�N�/����?�1�0�B���3�A�"�N�P�-��/�.�.�� �"��Qϊ0�-�D�o�  �&����#�]�M�#.�O������"�$��/����N�=�]���1��
���_�M�. �.�=�͊a�#�P��&/4�n����#� �1��"��@� ���@� !�2/=�� ��1� � ��N��C�����,#�Q����1��$���,4��$0�1 ��� �2�`����.�3>�@ �� �3�. ��Q�Q�O��/�4�!�3��.�+��o�2��$���j
�S���Q�!����E�$f� �0� �-��  3��;��4��4�;�#�5��`���A�"��%1��E�찊;�B�@��C#-����2���.#��E��l�<�>
�C5N�p;��=��!��!��B���3�#�֤_�2$��4���6��O���1����	�c�.И#�V�-����$,�D�Ҕ_���dˤ�@��/�3�#���S��.�U� �C�� ����4�/��1�V:�`ِ��.�/�B��?����L�?�4���U��D����Nϔ3�GM�A�3��^�+�7�>���� �����2���A��A��R��A�B��2�-��'��@�B�0�  ���T���ބT���m��� �Aݔ�m��4���B��0�R��#M�! Rݤ�@�F-�,�l�@���� ܤ!�$��A��?���1���4��P�V+��4�!�� ��4���b��o� �d��"�!#?�4��1*�,�� �c�=����N���j�b�����?����� 3�C!���#��"��0��B����O�#���M�!%,�P��"1�&M�"��A��R��,� 2>��-�N ����K�3,�0��s��bѤA�1�����3��3є/��C�>Ҙ��4,��A�.�U���T��>���?�A��GL�d�"��?��!�2��/�`�0ک�_�D ��C��V���>�� �_���M����ڤ �4/����.�N�E��R��Q�[�S�C�]�/�N�A�!�"                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                ��������������������������������                                �������������������������������� Z K � P d d d d d � � � � � d d��������������������������� U � � � 0 � � v P � � P P P P � ���������������������PP��                                ���$�$�	���c   a 8 � � � �               ��������   4 , d d j �             V   ����� ���@�@�@�@��        �� ; 4 ; / J C 4 E YD # � 3 & { �� � � � � � � � � �� ��� ��� �                 B            ������[�mX�X�X�X�������������~ �� � � �� ���  � �   ����8�                                                            ��������������������������������  ��  ��          4 ��  � F     �
�
��P!:Y	�1��	 
�j5�����������������������������������������������������������������               ��������������������� �����  &\%      �K    ��   ��������%����������4��                  >      &>    ��>������&>�������3�������7�������������                       ����������������������������������� �������x����/����~������� ����~���� �����]��  �� P��Z                                 �"�FV  �"�FV   K�FV                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        